#
#   VizieR Astronomical Server vizier.u-strasbg.fr
#    Date: 2017-08-24T13:58:22 [V1.99+ (14-Oct-2013)]
#   In case of problem, please report to:	cds-question@unistra.fr
#
#
#Coosys	J2000:	eq_FK5 J2000
#INFO	votable-version=1.99+ (14-Oct-2013)	
#INFO	-ref=VIZ599eafbf9987	
#INFO	-out.max=99999	
#INFO	queryParameters=16	
#-oc.form=dec
#-out.max=99999
#-out.all=2
#-order=I
#-nav=cat:J/ApJ/829/93&tab:{J/ApJ/829/93/table2}&key:source=J/ApJ/829/93/table2&HTTPPRM:&&-ref=VIZ599eafbf9987&-out.max=99999&-out.form=HTML Table&-out.all=2&-order=I&-oc.form=sexa&-out.src=J/ApJ/829/93/table2&-out=ID&-out=Line&-out=f_Line&-out=Flux&-out=b_Flux&-out=B_Flux&-out=UpLim&-meta.ucd=2&-meta=1&-meta.foot=1&-usenav=1&-bmark=POST&
#-order=I
#-source= J/ApJ/829/93/table2
#-order=I
#-out.src=J/ApJ/829/93/table2
#-out=ID
#-out=Line
#-out=f_Line
#-out=Flux
#-out=b_Flux
#-out=B_Flux
#-out=UpLim
#

#RESOURCE=yCat_18290093
#Name: J/ApJ/829/93
#Title: CO, [CI] and [NII] lines from Herschel spectra (Kamenetzky+, 2016)
#Table	J_ApJ_829_93_table2:
#Name: J/ApJ/829/93/table2
#Title: Line fluxes and uncertainty ranges from SPIRE FTS
#Column	ID	(a16)	Galaxy identifier \linkRole{observations data (table 1)}	[ucd=meta.id;meta.main]
#Column	Line	(A7)	Line identifier	[ucd=meta.id;spect.line]
#Column	f_Line	(A1)	[X] Line is resolved?	[ucd=meta.code]
#Column	Flux	(E8.1)	[14/89800] Median line flux in Line	[ucd=phot.flux.density;stat.median]
#Column	b_Flux	(E8.1)	Lower 1{sigma} boundary for Flux	[ucd=phot.flux.density;stat.min]
#Column	B_Flux	(E8.1)	Upper 1{sigma} boundary for Flux	[ucd=phot.flux.density;stat.max]
#Column	UpLim	(E8.1)	? The 3{sigma} upper limit on the Line flux (1)	[ucd=phot.flux.density;stat.max]
ID|Line|f_Line|Flux|b_Flux|B_Flux|UpLim
 | | |Jy.km/s|Jy.km/s|Jy.km/s|Jy.km/s
----------------|-------|-|--------|--------|--------|--------
NGC0023         |CI1-0  | | 2.6e+02| 6.8e+01| 5.6e+02| 8.0e+02
NGC0023         |CI2-1  | | 3.8e+02| 3.1e+02| 4.6e+02|
NGC0023         |CO4-3  | | 3.1e+02| 7.2e+01| 6.1e+02| 1.2e+03
NGC0023         |CO5-4  | | 7.4e+02| 5.8e+02| 9.7e+02|
NGC0023         |CO6-5  | | 4.2e+02| 3.3e+02| 4.9e+02|
NGC0023         |CO7-6  | | 3.2e+02| 2.4e+02| 4.0e+02|
NGC0023         |CO8-7  | | 2.5e+02| 1.2e+02| 3.8e+02| 5.7e+02
NGC0023         |CO9-8  | | 1.2e+02| 2.5e+01| 2.9e+02| 5.6e+02
NGC0023         |CO10-9 | | 2.2e+02| 5.5e+01| 3.6e+02| 5.3e+02
NGC0023         |CO12-11| | 7.8e+01| 1.8e+01| 1.9e+02| 3.3e+02
NGC0023         |CO13-12| | 2.3e+02| 9.7e+01| 3.6e+02| 4.8e+02
NGC0023         |NII    |X| 2.6e+03| 2.5e+03| 2.8e+03|
NGC34           |CI1-0  | | 5.0e+02| 3.4e+02| 6.4e+02|
NGC34           |CI2-1  | | 4.3e+02| 3.8e+02| 4.7e+02|
NGC34           |CO5-4  | | 7.9e+02| 6.9e+02| 8.8e+02|
NGC34           |CO6-5  | | 9.7e+02| 9.1e+02| 1.0e+03|
NGC34           |CO7-6  | | 9.5e+02| 9.1e+02| 9.9e+02|
NGC34           |CO8-7  | | 8.6e+02| 7.8e+02| 9.2e+02|
NGC34           |CO9-8  | | 6.2e+02| 5.7e+02| 6.7e+02|
NGC34           |CO10-9 | | 4.6e+02| 4.2e+02| 5.0e+02|
NGC34           |CO11-10| | 4.0e+02| 3.6e+02| 4.4e+02|
NGC34           |CO12-11| | 2.7e+02| 2.4e+02| 3.0e+02|
NGC34           |CO13-12| | 2.0e+02| 1.6e+02| 2.4e+02|
NGC34           |NII    |X| 7.1e+02| 6.6e+02| 7.6e+02|
MCG-02-01-051   |CI1-0  | | 1.1e+02| 3.2e+01| 2.2e+02| 3.9e+02
MCG-02-01-051   |CI2-1  | | 2.2e+02| 1.7e+02| 2.7e+02|
MCG-02-01-051   |CO5-4  | | 3.2e+02| 2.0e+02| 4.4e+02|
MCG-02-01-051   |CO6-5  | | 3.9e+02| 3.2e+02| 4.5e+02|
MCG-02-01-051   |CO7-6  | | 2.4e+02| 1.9e+02| 2.9e+02|
MCG-02-01-051   |CO8-7  | | 2.0e+02| 1.2e+02| 2.7e+02|
MCG-02-01-051   |CO9-8  | | 2.6e+02| 1.7e+02| 3.7e+02|
MCG-02-01-051   |CO10-9 | | 1.7e+02| 9.2e+01| 2.3e+02|
MCG-02-01-051   |CO11-10| | 3.3e+01| 5.4e+00| 7.5e+01| 1.4e+02
MCG-02-01-051   |CO12-11| | 1.1e+02| 5.3e+01| 1.7e+02| 2.4e+02
MCG-02-01-051   |CO13-12| | 7.1e+01| 1.9e+01| 1.2e+02| 2.2e+02
MCG-02-01-051   |NII    | | 5.6e+02| 5.1e+02| 6.1e+02|
IC10-B11-1      |CI1-0  | | 2.4e+02| 1.4e+02| 3.2e+02| 4.4e+02
IC10-B11-1      |CI2-1  | | 5.9e+02| 5.4e+02| 6.4e+02|
IC10-B11-1      |CO4-3  | | 6.6e+02| 5.5e+02| 7.6e+02|
IC10-B11-1      |CO5-4  | | 8.2e+02| 7.3e+02| 9.0e+02|
IC10-B11-1      |CO6-5  | | 7.8e+02| 7.2e+02| 8.2e+02|
IC10-B11-1      |CO7-6  | | 5.9e+02| 5.4e+02| 6.5e+02|
IC10-B11-1      |CO8-7  | | 3.2e+02| 2.3e+02| 3.9e+02|
IC10-B11-1      |CO9-8  | | 3.0e+02| 1.7e+02| 4.2e+02|
IC10-B11-1      |CO10-9 | | 2.0e+02| 9.8e+01| 2.8e+02| 4.6e+02
IC10-B11-1      |CO11-10| | 1.3e+02| 4.2e+01| 2.3e+02| 4.1e+02
IC10-B11-1      |CO12-11| | 1.3e+02| 5.1e+01| 2.2e+02| 3.5e+02
IC10-B11-1      |CO13-12| | 1.3e+02| 4.6e+01| 2.4e+02| 3.7e+02
IC10-B11-1      |NII    | | 1.6e+03| 1.5e+03| 1.8e+03|
IRAS 00188-0856 |CI2-1  | | 9.2e+01| 4.0e+01| 1.3e+02|
IRAS 00188-0856 |CO5-4  | | 6.7e+01| 1.1e+01| 1.8e+02| 3.4e+02
IRAS 00188-0856 |CO6-5  | | 4.0e+01| 5.7e+00| 9.9e+01| 2.0e+02
IRAS 00188-0856 |CO7-6  | | 1.1e+02| 6.6e+01| 1.5e+02|
IRAS 00188-0856 |CO8-7  | | 1.0e+02| 7.2e+01| 1.4e+02|
IRAS 00188-0856 |CO10-9 | | 9.2e+01| 4.3e+01| 1.3e+02| 2.1e+02
IRAS 00188-0856 |CO11-10| | 2.8e+01| 5.8e+00| 6.6e+01| 1.1e+02
IRAS 00188-0856 |CO12-11| | 7.3e+01| 4.1e+01| 1.1e+02| 1.6e+02
IRAS 00188-0856 |NII    | | 8.6e+01| 5.4e+01| 1.2e+02|
ESO350-IG038    |CI2-1  | | 1.0e+02| 3.5e+01| 1.9e+02| 3.0e+02
ESO350-IG038    |CO5-4  | | 5.0e+01| 3.9e-01| 1.4e+02| 3.4e+02
ESO350-IG038    |CO7-6  | | 1.2e+02| 4.2e+01| 2.1e+02| 3.1e+02
ESO350-IG038    |CO9-8  | | 1.2e+02| 2.7e+01| 2.9e+02| 5.0e+02
ESO350-IG038    |CO10-9 | | 8.2e+01| 1.1e+01| 2.1e+02| 4.2e+02
ESO350-IG038    |CO11-10| | 1.2e+02| 2.6e+01| 2.1e+02| 3.3e+02
ESO350-IG038    |CO12-11| | 4.2e+01| 5.4e+00| 1.0e+02| 1.9e+02
ESO350-IG038    |CO13-12| | 5.1e+01| 8.7e+00| 1.2e+02| 2.8e+02
ESO350-IG038    |NII    | | 4.8e+02| 3.8e+02| 5.8e+02|
NGC205-copeak   |CI1-0  | | 2.2e+02| 1.1e+02| 3.5e+02| 4.9e+02
NGC205-copeak   |CI2-1  | | 1.5e+01| 2.4e+00| 4.0e+01| 8.4e+01
NGC205-copeak   |CO4-3  | | 2.4e+02| 1.0e+02| 3.5e+02| 5.5e+02
NGC205-copeak   |CO6-5  | | 3.4e+01| 6.9e+00| 7.6e+01| 1.2e+02
NGC205-copeak   |CO7-6  | | 3.4e+01| 1.4e+01| 5.9e+01| 1.1e+02
NGC205-copeak   |CO8-7  | | 9.3e+01| 4.7e+01| 1.5e+02| 2.2e+02
NGC205-copeak   |CO9-8  | | 7.9e+01| 2.4e+01| 1.8e+02| 3.3e+02
NGC205-copeak   |CO10-9 | | 6.8e+01| 1.1e+01| 1.4e+02| 2.4e+02
NGC205-copeak   |CO11-10| | 1.6e+02| 8.5e+01| 2.4e+02| 3.5e+02
NGC205-copeak   |CO13-12| | 2.0e+02| 1.3e+02| 2.7e+02|
IRAS 00397-1312 |CI2-1  | | 5.1e+01| 1.5e+01| 9.4e+01| 1.6e+02
IRAS 00397-1312 |CO5-4  | | 2.2e+02| 6.6e+01| 3.4e+02| 5.5e+02
IRAS 00397-1312 |CO6-5  | | 1.1e+02| 3.1e+01| 2.0e+02| 3.6e+02
IRAS 00397-1312 |CO8-7  | | 6.4e+01| 2.7e+01| 9.9e+01| 1.6e+02
IRAS 00397-1312 |CO12-11| | 9.0e+01| 5.2e+01| 1.3e+02| 1.8e+02
IRAS 00397-1312 |CO13-12| | 4.0e+01| 1.1e+01| 7.3e+01| 1.2e+02
IRAS 00397-1312 |NII    | | 4.7e+01| 1.6e+01| 7.4e+01| 1.2e+02
NGC0232a        |CI1-0  | | 7.9e+02| 4.5e+02| 1.3e+03|
NGC0232a        |CI2-1  | | 8.1e+02| 7.4e+02| 8.8e+02|
NGC0232a        |CO5-4  | | 1.0e+03| 8.4e+02| 1.3e+03|
NGC0232a        |CO6-5  | | 8.3e+02| 7.3e+02| 9.3e+02|
NGC0232a        |CO7-6  | | 6.3e+02| 5.6e+02| 7.0e+02|
NGC0232a        |CO8-7  | | 4.6e+02| 3.7e+02| 5.4e+02|
NGC0232a        |CO9-8  | | 2.0e+02| 1.1e+02| 3.2e+02| 5.0e+02
NGC0232a        |CO10-9 | | 2.4e+02| 1.6e+02| 3.3e+02|
NGC0232a        |CO11-10| | 7.2e+01| 1.9e+01| 1.6e+02| 2.9e+02
NGC0232a        |CO12-11| | 5.0e+01| 8.9e+00| 1.0e+02| 1.8e+02
NGC0232a        |CO13-12| | 8.2e+01| 2.8e+01| 1.4e+02| 2.6e+02
NGC0232a        |NII    |X| 2.2e+03| 2.1e+03| 2.2e+03|
NGC253          |CI1-0  | | 2.6e+04| 2.5e+04| 2.7e+04|
NGC253          |CI2-1  | | 4.0e+04| 3.9e+04| 4.1e+04|
NGC253          |CO4-3  | | 7.5e+04| 7.4e+04| 7.7e+04|
NGC253          |CO5-4  | | 8.4e+04| 8.4e+04| 8.5e+04|
NGC253          |CO6-5  | | 7.4e+04| 7.4e+04| 7.5e+04|
NGC253          |CO7-6  | | 6.3e+04| 6.2e+04| 6.4e+04|
NGC253          |CO8-7  | | 5.2e+04| 5.0e+04| 5.3e+04|
NGC253          |CO9-8  | | 4.2e+04| 4.0e+04| 4.4e+04|
NGC253          |CO10-9 | | 3.0e+04| 2.8e+04| 3.1e+04|
NGC253          |CO11-10| | 2.2e+04| 2.0e+04| 2.4e+04|
NGC253          |CO12-11| | 1.6e+04| 1.5e+04| 1.7e+04|
NGC253          |CO13-12| | 8.9e+03| 6.4e+03| 1.2e+04| 1.8e+04
NGC253          |NII    | | 3.6e+04| 3.4e+04| 3.8e+04|
I Zw 1          |CI1-0  | | 2.3e+02| 8.0e+01| 5.1e+02| 7.1e+02
I Zw 1          |CI2-1  | | 9.4e+01| 5.4e+01| 1.4e+02| 2.0e+02
I Zw 1          |CO6-5  | | 7.3e+01| 2.3e+01| 1.3e+02| 2.3e+02
I Zw 1          |CO7-6  | | 5.7e+01| 1.8e+01| 9.8e+01| 1.7e+02
I Zw 1          |CO8-7  | | 8.7e+01| 3.2e+01| 1.3e+02| 2.0e+02
I Zw 1          |CO9-8  | | 2.1e+02| 1.4e+02| 2.8e+02|
I Zw 1          |CO10-9 | | 4.1e+01| 9.6e+00| 8.8e+01| 1.6e+02
I Zw 1          |CO11-10| | 5.0e+01| 1.9e+01| 9.8e+01| 1.6e+02
I Zw 1          |CO12-11| | 1.7e+01| 2.2e+00| 4.2e+01| 1.0e+02
I Zw 1          |CO13-12| | 3.0e+01| 8.5e+00| 6.2e+01| 1.3e+02
I Zw 1          |NII    | | 2.3e+02| 1.9e+02| 2.7e+02|
MCG+12-02-001   |CI1-0  | | 4.4e+02| 3.0e+02| 5.6e+02|
MCG+12-02-001   |CI2-1  | | 6.3e+02| 6.0e+02| 6.7e+02|
MCG+12-02-001   |CO4-3  | | 1.2e+03| 1.1e+03| 1.4e+03|
MCG+12-02-001   |CO5-4  | | 1.2e+03| 1.1e+03| 1.3e+03|
MCG+12-02-001   |CO6-5  | | 9.5e+02| 9.1e+02| 9.8e+02|
MCG+12-02-001   |CO7-6  | | 6.5e+02| 6.2e+02| 6.9e+02|
MCG+12-02-001   |CO8-7  | | 5.2e+02| 4.5e+02| 5.7e+02|
MCG+12-02-001   |CO9-8  | | 4.6e+02| 4.0e+02| 5.2e+02|
MCG+12-02-001   |CO10-9 | | 2.7e+02| 2.2e+02| 3.2e+02|
MCG+12-02-001   |CO11-10| | 2.9e+02| 2.4e+02| 3.4e+02|
MCG+12-02-001   |CO12-11| | 8.3e+01| 3.8e+01| 1.2e+02| 1.9e+02
MCG+12-02-001   |CO13-12| | 9.4e+01| 3.1e+01| 1.7e+02| 2.6e+02
MCG+12-02-001   |NII    | | 1.8e+03| 1.7e+03| 1.8e+03|
NGC0317B        |CI1-0  | | 1.6e+02| 6.0e+01| 2.6e+02| 4.3e+02
NGC0317B        |CI2-1  | | 4.3e+02| 3.8e+02| 4.7e+02|
NGC0317B        |CO4-3  | | 1.6e+02| 4.4e+01| 2.5e+02| 4.1e+02
NGC0317B        |CO5-4  | | 4.2e+02| 3.5e+02| 5.1e+02|
NGC0317B        |CO6-5  | | 3.6e+02| 3.1e+02| 4.1e+02|
NGC0317B        |CO7-6  | | 3.8e+02| 3.3e+02| 4.2e+02|
NGC0317B        |CO8-7  | | 1.9e+02| 1.4e+02| 2.5e+02|
NGC0317B        |CO9-8  | | 3.3e+02| 2.4e+02| 4.1e+02|
NGC0317B        |CO10-9 | | 1.2e+02| 5.5e+01| 2.0e+02| 3.0e+02
NGC0317B        |CO11-10| | 2.6e+02| 2.0e+02| 3.3e+02|
NGC0317B        |CO13-12| | 5.6e+01| 1.9e+01| 1.0e+02| 1.8e+02
NGC0317B        |NII    | | 6.4e+02| 5.8e+02| 7.0e+02|
IRAS 01003-2238 |CI2-1  | | 6.8e+01| 3.1e+01| 9.7e+01| 1.5e+02
IRAS 01003-2238 |CO6-5  | | 7.8e+01| 2.4e+01| 1.6e+02| 2.3e+02
IRAS 01003-2238 |CO7-6  | | 4.6e+01| 2.1e+01| 7.5e+01| 1.2e+02
IRAS 01003-2238 |CO8-7  | | 4.0e+01| 9.8e+00| 7.6e+01| 1.1e+02
IRAS 01003-2238 |CO10-9 | | 1.3e+02| 7.6e+01| 1.8e+02|
IRAS 01003-2238 |CO11-10| | 8.3e+01| 4.8e+01| 1.1e+02| 1.7e+02
IRAS 01003-2238 |CO12-11| | 4.9e+01| 1.5e+01| 9.9e+01| 1.4e+02
IRAS 01003-2238 |CO13-12| | 3.6e+01| 1.1e+01| 6.5e+01| 9.9e+01
3C 31           |CI1-0  | | 5.6e+01| 1.1e+01| 1.2e+02| 2.3e+02
3C 31           |CI2-1  | | 3.2e+01| 1.3e+01| 4.7e+01| 7.4e+01
3C 31           |CO4-3  | | 1.4e+02| 4.2e+01| 2.4e+02| 4.3e+02
3C 31           |CO6-5  | | 2.7e+01| 7.5e+00| 5.2e+01| 8.8e+01
3C 31           |CO7-6  | | 3.8e+01| 2.2e+01| 5.2e+01|
3C 31           |CO10-9 | | 7.0e+01| 3.7e+01| 1.0e+02|
3C 31           |CO12-11| | 5.0e+01| 2.2e+01| 7.5e+01| 1.2e+02
3C 31           |NII    | | 8.3e+01| 5.6e+01| 1.1e+02|
IC1623          |CI1-0  | | 1.8e+03| 1.4e+03| 2.1e+03|
IC1623          |CI2-1  | | 1.4e+03| 1.3e+03| 1.4e+03|
IC1623          |CO5-4  | | 3.4e+03| 3.2e+03| 3.5e+03|
IC1623          |CO6-5  | | 1.9e+03| 1.8e+03| 2.0e+03|
IC1623          |CO7-6  | | 1.2e+03| 1.2e+03| 1.3e+03|
IC1623          |CO8-7  | | 8.2e+02| 7.5e+02| 8.8e+02|
IC1623          |CO9-8  | | 5.6e+02| 4.6e+02| 6.4e+02|
IC1623          |CO10-9 | | 3.1e+02| 2.5e+02| 3.9e+02|
IC1623          |CO11-10| | 1.5e+02| 7.4e+01| 2.3e+02| 3.7e+02
IC1623          |CO12-11| | 2.0e+02| 1.4e+02| 2.7e+02|
IC1623          |CO13-12| | 2.6e+02| 1.6e+02| 3.4e+02|
IC1623          |NII    |X| 3.0e+03| 2.9e+03| 3.1e+03|
MCG-03-04-014   |CI1-0  | | 4.0e+02| 2.0e+02| 5.8e+02| 1.0e+03
MCG-03-04-014   |CI2-1  | | 3.8e+02| 3.1e+02| 4.1e+02|
MCG-03-04-014   |CO5-4  | | 5.3e+02| 3.9e+02| 7.0e+02|
MCG-03-04-014   |CO6-5  | | 5.1e+02| 4.5e+02| 5.7e+02|
MCG-03-04-014   |CO7-6  | | 3.9e+02| 3.4e+02| 4.5e+02|
MCG-03-04-014   |CO8-7  | | 1.6e+02| 8.2e+01| 2.4e+02|
MCG-03-04-014   |CO9-8  | | 9.0e+01| 2.2e+01| 1.4e+02| 2.5e+02
MCG-03-04-014   |CO10-9 | | 6.9e+01| 2.8e+01| 1.2e+02| 1.9e+02
MCG-03-04-014   |CO11-10| | 5.1e+01| 1.8e+01| 9.5e+01| 1.4e+02
MCG-03-04-014   |CO12-11| | 8.2e+01| 3.7e+01| 1.3e+02| 2.1e+02
MCG-03-04-014   |CO13-12| | 7.9e+01| 3.1e+01| 1.3e+02| 1.8e+02
MCG-03-04-014   |NII    |X| 1.8e+03| 1.8e+03| 1.9e+03|
ESO244-G012     |CI2-1  | | 4.3e+02| 3.6e+02| 5.2e+02|
ESO244-G012     |CO5-4  | | 4.7e+02| 2.3e+02| 6.6e+02| 9.5e+02
ESO244-G012     |CO6-5  | | 8.9e+02| 7.7e+02| 1.0e+03|
ESO244-G012     |CO7-6  | | 3.8e+02| 3.1e+02| 4.6e+02|
ESO244-G012     |CO8-7  | | 3.4e+02| 2.4e+02| 4.3e+02|
ESO244-G012     |CO9-8  | | 1.8e+02| 7.7e+01| 3.2e+02| 4.8e+02
ESO244-G012     |CO10-9 | | 1.9e+02| 9.5e+01| 2.8e+02| 3.9e+02
ESO244-G012     |CO11-10| | 1.5e+02| 5.6e+01| 2.3e+02| 3.5e+02
ESO244-G012     |CO12-11| | 1.1e+02| 3.4e+01| 1.8e+02| 3.1e+02
ESO244-G012     |CO13-12| | 1.1e+02| 3.6e+01| 1.9e+02| 3.1e+02
ESO244-G012     |NII    | | 6.0e+02| 5.3e+02| 6.7e+02|
CGCG436-030     |CI1-0  | | 3.8e+02| 1.5e+02| 6.2e+02| 9.6e+02
CGCG436-030     |CI2-1  | | 3.4e+02| 2.9e+02| 4.0e+02|
CGCG436-030     |CO5-4  | | 6.1e+02| 4.8e+02| 7.9e+02|
CGCG436-030     |CO6-5  | | 5.3e+02| 4.6e+02| 6.0e+02|
CGCG436-030     |CO7-6  | | 4.3e+02| 3.8e+02| 5.0e+02|
CGCG436-030     |CO8-7  | | 4.5e+02| 3.8e+02| 5.2e+02|
CGCG436-030     |CO9-8  | | 1.9e+02| 1.2e+02| 2.8e+02|
CGCG436-030     |CO10-9 | | 1.5e+02| 8.3e+01| 2.0e+02|
CGCG436-030     |CO11-10| | 2.2e+02| 1.6e+02| 2.8e+02|
CGCG436-030     |CO12-11| | 4.7e+01| 1.4e+01| 9.0e+01| 1.6e+02
CGCG436-030     |CO13-12| | 5.6e+01| 1.7e+01| 1.0e+02| 1.7e+02
CGCG436-030     |NII    | | 3.8e+02| 3.4e+02| 4.3e+02|
ESO353-G020     |CI1-0  | | 3.2e+02| 1.2e+02| 6.0e+02| 9.6e+02
ESO353-G020     |CI2-1  | | 8.3e+02| 7.8e+02| 8.9e+02|
ESO353-G020     |CO4-3  | | 5.8e+02| 3.5e+02| 8.4e+02|
ESO353-G020     |CO5-4  | | 1.1e+03| 9.3e+02| 1.2e+03|
ESO353-G020     |CO6-5  | | 7.4e+02| 6.7e+02| 8.1e+02|
ESO353-G020     |CO7-6  | | 5.6e+02| 4.8e+02| 6.2e+02|
ESO353-G020     |CO8-7  | | 1.9e+02| 1.2e+02| 2.8e+02|
ESO353-G020     |CO9-8  | | 6.4e+01| 1.2e+01| 1.4e+02| 2.8e+02
ESO353-G020     |CO10-9 | | 9.4e+01| 3.5e+01| 1.8e+02| 2.7e+02
ESO353-G020     |CO11-10| | 1.3e+02| 5.4e+01| 2.0e+02| 3.3e+02
ESO353-G020     |CO12-11| | 1.1e+02| 4.4e+01| 1.9e+02| 2.8e+02
ESO353-G020     |NII    |X| 3.4e+03| 3.3e+03| 3.5e+03|
IIIZw035             |CI1-0   |        |  1.66e+02|  7.23e+01|  2.57e+02|  3.85e+02 
IIIZw035             |CI2-1   |        |  1.63e+02|  1.27e+02|  1.90e+02|           
IIIZw035             |CO5-4   |        |  1.21e+02|  5.45e+01|  2.09e+02|  3.36e+02
IIIZw035             |CO6-5   |        |  2.42e+02|  1.95e+02|  2.86e+02|           
IIIZw035             |CO7-6   |        |  3.05e+02|  2.69e+02|  3.39e+02|           
IIIZw035             |CO8-7   |        |  3.68e+02|  3.22e+02|  4.16e+02|           
IIIZw035             |CO9-8   |        |  3.52e+02|  2.55e+02|  4.45e+02|           
IIIZw035             |CO10-9  |        |  4.23e+02|  3.60e+02|  4.93e+02|           
IIIZw035             |CO11-10 |        |  1.50e+02|  8.86e+01|  2.03e+02|  3.09e+02 
IIIZw035             |CO12-11 |        |  1.58e+02|  9.95e+01|  2.18e+02|           
IIIZw035             |CO13-12 |        |  8.08e+01|  3.49e+01|  1.24e+02|  2.31e+02 
IIIZw035             |NII     |        |  9.04e+01|  3.84e+01|  1.40e+02|  2.20e+02
NGC0695         |CI1-0  | | 5.8e+02| 2.1e+02| 9.0e+02| 1.4e+03
NGC0695         |CI2-1  | | 4.7e+02| 4.2e+02| 5.3e+02|
NGC0695         |CO5-4  | | 1.1e+03| 8.9e+02| 1.3e+03|
NGC0695         |CO6-5  | | 4.7e+02| 3.7e+02| 5.6e+02|
NGC0695         |CO7-6  | | 3.7e+02| 3.2e+02| 4.3e+02|
NGC0695         |CO8-7  | | 2.3e+02| 1.6e+02| 2.9e+02|
NGC0695         |CO9-8  | | 1.1e+02| 4.2e+01| 2.1e+02| 3.8e+02
NGC0695         |CO10-9 | | 4.0e+01| 6.1e+00| 9.2e+01| 1.5e+02
NGC0695         |CO11-10| | 3.7e+01| 6.0e+00| 9.0e+01| 1.5e+02
NGC0695         |CO13-12| | 5.4e+01| 1.4e+01| 1.0e+02| 1.7e+02
NGC0695         |NII    | | 2.4e+03| 2.3e+03| 2.4e+03|
Mrk 1014        |CI2-1  | | 9.6e+01| 4.9e+01| 1.5e+02| 2.4e+02
Mrk 1014        |CO5-4  | | 3.2e+02| 1.5e+02| 4.7e+02| 6.3e+02
Mrk 1014        |CO6-5  | | 1.4e+02| 4.5e+01| 2.5e+02| 3.5e+02
Mrk 1014        |CO7-6  | | 8.1e+01| 3.7e+01| 1.4e+02| 2.4e+02
Mrk 1014        |CO10-9 | | 3.5e+01| 7.7e+00| 6.5e+01| 1.0e+02
Mrk 1014        |CO11-10| | 2.4e+01| 7.5e+00| 5.6e+01| 8.7e+01
Mrk 1014        |CO13-12| | 3.7e+01| 1.3e+01| 6.7e+01| 1.2e+02
Mrk 1014        |NII    | | 9.5e+01| 6.3e+01| 1.2e+02|
NGC0828         |CI1-0  | | 7.0e+02| 4.4e+02| 1.0e+03| 1.5e+03
NGC0828         |CI2-1  | | 6.2e+02| 5.4e+02| 7.0e+02|
NGC0828         |CO4-3  | | 9.3e+02| 6.0e+02| 1.3e+03| 1.9e+03
NGC0828         |CO5-4  | | 7.6e+02| 5.3e+02| 1.0e+03|
NGC0828         |CO6-5  | | 8.2e+02| 6.8e+02| 9.4e+02|
NGC0828         |CO7-6  | | 1.6e+02| 7.4e+01| 2.4e+02| 3.5e+02
NGC0828         |CO8-7  | | 1.7e+02| 6.2e+01| 3.0e+02| 5.3e+02
NGC0828         |CO10-9 | | 1.8e+02| 6.5e+01| 3.0e+02| 5.0e+02
NGC0828         |CO11-10| | 9.7e+01| 2.9e+01| 2.0e+02| 3.6e+02
NGC0828         |CO12-11| | 1.2e+02| 3.7e+01| 2.0e+02| 3.8e+02
NGC0828         |NII    |X| 7.2e+03| 7.0e+03| 7.4e+03|
NGC0877a        |CI1-0  | | 3.6e+02| 1.6e+02| 5.8e+02| 8.6e+02
NGC0877a        |CI2-1  | | 3.9e+02| 3.0e+02| 4.8e+02|
NGC0877a        |CO4-3  | | 3.7e+02| 1.6e+02| 6.3e+02| 8.9e+02
NGC0877a        |CO5-4  | | 2.9e+02| 1.2e+02| 4.6e+02| 8.1e+02
NGC0877a        |CO6-5  | | 2.4e+02| 1.4e+02| 3.4e+02|
NGC0877a        |CO7-6  | | 2.2e+02| 1.3e+02| 3.1e+02|
NGC0877a        |CO8-7  | | 1.3e+02| 3.9e+01| 2.3e+02| 4.0e+02
NGC0877a        |CO9-8  | | 6.5e+02| 3.3e+02| 9.6e+02|
NGC0877a        |CO10-9 | | 1.5e+02| 2.4e+01| 4.0e+02| 6.5e+02
NGC0877a        |CO11-10| | 4.6e+02| 2.3e+02| 6.9e+02| 1.1e+03
NGC0877a        |CO13-12| | 5.4e+02| 2.2e+02| 8.0e+02| 1.2e+03
NGC0877a        |NII    | | 4.5e+03| 4.2e+03| 4.7e+03|
NGC891-1        |CI1-0  | | 2.2e+03| 1.9e+03| 2.5e+03|
NGC891-1        |CI2-1  | | 1.8e+03| 1.7e+03| 2.0e+03|
NGC891-1        |CO4-3  | | 2.2e+03| 1.9e+03| 2.6e+03|
NGC891-1        |CO5-4  | | 2.0e+03| 1.6e+03| 2.3e+03|
NGC891-1        |CO6-5  | | 1.3e+03| 1.1e+03| 1.4e+03|
NGC891-1        |CO7-6  | | 7.8e+02| 6.4e+02| 9.2e+02|
NGC891-1        |CO8-7  | | 4.8e+02| 2.3e+02| 7.4e+02| 9.6e+02
NGC891-1        |CO9-8  | | 1.9e+02| 3.0e+01| 4.2e+02| 8.2e+02
NGC891-1        |CO10-9 | | 4.3e+02| 1.9e+02| 7.1e+02| 1.5e+03
NGC891-1        |CO11-10| | 3.2e+02| 7.4e+01| 5.9e+02| 9.7e+02
NGC891-1        |CO12-11| | 1.4e+02| 1.6e+01| 3.1e+02| 5.6e+02
NGC891-1        |NII    | | 1.6e+04| 1.6e+04| 1.6e+04|
UGC01845        |CI1-0  | | 2.0e+02| 3.8e+01| 3.6e+02| 6.4e+02
UGC01845        |CI2-1  | | 3.9e+02| 3.2e+02| 4.5e+02|
UGC01845        |CO4-3  | | 1.3e+02| 1.4e+01| 3.4e+02| 8.2e+02
UGC01845        |CO5-4  | | 6.5e+02| 5.1e+02| 8.0e+02|
UGC01845        |CO6-5  | | 4.6e+02| 3.9e+02| 5.4e+02|
UGC01845        |CO7-6  | | 3.7e+02| 3.0e+02| 4.3e+02|
UGC01845        |CO8-7  | | 2.4e+02| 1.4e+02| 3.3e+02| 4.6e+02
UGC01845        |CO9-8  | | 1.5e+02| 4.9e+01| 2.8e+02| 4.8e+02
UGC01845        |CO10-9 | | 1.8e+02| 5.9e+01| 2.8e+02| 4.1e+02
UGC01845        |CO12-11| | 1.1e+02| 3.4e+01| 2.0e+02| 3.4e+02
UGC01845        |CO13-12| | 7.7e+01| 2.1e+01| 1.4e+02| 2.7e+02
UGC01845        |NII    |X| 2.8e+03| 2.6e+03| 2.9e+03|
NGC0958         |CI1-0  | | 2.0e+02| 7.2e+01| 3.5e+02| 5.2e+02
NGC0958         |CI2-1  | | 1.3e+02| 7.1e+01| 2.0e+02|
NGC0958         |CO5-4  | | 4.1e+01| 1.9e+00| 1.2e+02| 2.7e+02
NGC0958         |CO6-5  | | 1.7e+02| 6.8e+01| 2.5e+02| 3.9e+02
NGC0958         |CO7-6  | | 8.2e+01| 2.8e+01| 1.4e+02| 2.2e+02
NGC0958         |CO9-8  | | 4.6e+02| 2.6e+02| 6.3e+02|
NGC0958         |CO10-9 | | 1.4e+02| 3.7e+01| 2.8e+02| 4.5e+02
NGC0958         |CO12-11| | 1.1e+02| 2.2e+01| 2.6e+02| 5.3e+02
NGC0958         |CO13-12| | 1.6e+02| 4.4e+01| 3.4e+02| 5.3e+02
NGC0958         |NII    |X| 3.6e+03| 3.3e+03| 3.8e+03|
0235+164        |CO8-7  | | 3.0e+01| 4.4e+00| 7.9e+01| 1.3e+02
NGC1068         |CI1-0  | | 8.6e+03| 8.1e+03| 8.9e+03|
NGC1068         |CI2-1  | | 1.1e+04| 1.1e+04| 1.1e+04|
NGC1068         |CO4-3  | | 1.4e+04| 1.3e+04| 1.4e+04|
NGC1068         |CO5-4  | | 1.2e+04| 1.2e+04| 1.2e+04|
NGC1068         |CO6-5  | | 1.1e+04| 1.1e+04| 1.1e+04|
NGC1068         |CO7-6  | | 7.5e+03| 7.3e+03| 7.8e+03|
NGC1068         |CO8-7  | | 6.4e+03| 5.8e+03| 6.8e+03|
NGC1068         |CO9-8  | | 7.6e+03| 7.0e+03| 8.2e+03|
NGC1068         |CO10-9 | | 7.0e+03| 6.5e+03| 7.4e+03|
NGC1068         |CO11-10| | 6.0e+03| 5.6e+03| 6.5e+03|
NGC1068         |CO12-11| | 5.3e+03| 4.9e+03| 5.7e+03|
NGC1068         |CO13-12| | 2.7e+03| 2.0e+03| 3.5e+03|
NGC1068         |NII    |X| 3.8e+04| 3.7e+04| 4.0e+04|
NGC1056         |CI1-0  | | 7.7e+01| 2.3e+01| 1.4e+02| 2.6e+02
NGC1056         |CI2-1  | | 2.4e+02| 1.8e+02| 2.9e+02|
NGC1056         |CO4-3  | | 6.5e+01| 1.6e+01| 1.2e+02| 2.1e+02
NGC1056         |CO5-4  | | 1.1e+02| 4.1e+01| 1.9e+02| 2.6e+02
NGC1056         |CO6-5  | | 1.7e+02| 1.2e+02| 2.2e+02|
NGC1056         |CO7-6  | | 1.7e+02| 1.2e+02| 2.2e+02|
NGC1056         |CO8-7  | | 1.0e+02| 3.8e+01| 1.8e+02| 3.1e+02
NGC1056         |CO9-8  | | 2.6e+02| 1.3e+02| 3.8e+02|
NGC1056         |CO10-9 | | 8.5e+01| 2.5e+01| 1.9e+02| 3.1e+02
NGC1056         |CO11-10| | 1.2e+02| 4.3e+01| 1.9e+02| 3.1e+02
NGC1056         |CO12-11| | 8.5e+01| 3.1e+01| 1.5e+02| 2.7e+02
NGC1056         |CO13-12| | 7.0e+01| 1.6e+01| 1.4e+02| 2.7e+02
NGC1056         |NII    | | 1.3e+03| 1.2e+03| 1.4e+03|
UGC02238        |CI1-0  | | 3.4e+02| 1.8e+02| 5.0e+02| 7.5e+02
UGC02238        |CI2-1  | | 4.0e+02| 3.6e+02| 4.4e+02|
UGC02238        |CO5-4  | | 5.0e+02| 4.2e+02| 5.9e+02|
UGC02238        |CO6-5  | | 3.4e+02| 2.9e+02| 4.0e+02|
UGC02238        |CO7-6  | | 1.6e+02| 1.2e+02| 2.1e+02|
UGC02238        |CO8-7  | | 7.5e+01| 2.4e+01| 1.4e+02| 2.8e+02
UGC02238        |CO9-8  | | 1.1e+02| 3.8e+01| 2.0e+02| 3.3e+02
UGC02238        |CO10-9 | | 1.0e+02| 3.4e+01| 1.7e+02| 3.0e+02
UGC02238        |CO11-10| | 8.1e+01| 2.7e+01| 1.7e+02| 3.3e+02
UGC02238        |NII    | | 2.2e+03| 2.2e+03| 2.3e+03|
NGC1097         |CI1-0  | | 2.5e+03| 2.2e+03| 2.8e+03|
NGC1097         |CI2-1  | | 2.5e+03| 2.4e+03| 2.6e+03|
NGC1097         |CO4-3  | | 3.6e+03| 3.2e+03| 3.9e+03|
NGC1097         |CO5-4  | | 3.4e+03| 3.2e+03| 3.7e+03|
NGC1097         |CO6-5  | | 2.7e+03| 2.6e+03| 2.8e+03|
NGC1097         |CO7-6  | | 1.6e+03| 1.5e+03| 1.7e+03|
NGC1097         |CO8-7  | | 6.4e+02| 4.3e+02| 8.1e+02|
NGC1097         |CO9-8  | | 4.4e+02| 1.8e+02| 6.4e+02| 9.0e+02
NGC1097         |CO10-9 | | 4.9e+02| 2.4e+02| 7.0e+02| 1.1e+03
NGC1097         |CO11-10| | 4.1e+02| 2.1e+02| 6.7e+02| 1.0e+03
NGC1097         |CO12-11| | 3.6e+02| 1.2e+02| 5.4e+02| 8.5e+02
NGC1097         |CO13-12| | 7.1e+02| 2.7e+02| 1.1e+03| 1.5e+03
NGC1097         |NII    |X| 1.9e+04| 1.8e+04| 1.9e+04|
UGC02369        |CI1-0  | | 9.0e+01| 2.4e+01| 1.6e+02| 3.0e+02
UGC02369        |CI2-1  | | 2.8e+02| 2.5e+02| 3.1e+02|
UGC02369        |CO5-4  | | 4.9e+02| 4.0e+02| 5.7e+02|
UGC02369        |CO6-5  | | 3.1e+02| 2.8e+02| 3.5e+02|
UGC02369        |CO7-6  | | 3.0e+02| 2.6e+02| 3.2e+02|
UGC02369        |CO8-7  | | 2.3e+02| 1.9e+02| 2.8e+02|
UGC02369        |CO9-8  | | 2.4e+02| 1.7e+02| 3.0e+02|
UGC02369        |CO10-9 | | 1.7e+02| 1.2e+02| 2.2e+02|
UGC02369        |CO12-11| | 7.6e+01| 1.4e+01| 1.2e+02| 1.8e+02
UGC02369        |CO13-12| | 9.8e+01| 3.4e+01| 1.4e+02| 2.1e+02
UGC02369        |NII    | | 8.6e+02| 8.1e+02| 9.1e+02|
NGC1222         |CI1-0  | | 2.4e+02| 1.3e+02| 3.4e+02|
NGC1222         |CI2-1  | | 2.2e+02| 1.9e+02| 2.5e+02|
NGC1222         |CO4-3  | | 2.6e+02| 1.4e+02| 3.8e+02|
NGC1222         |CO5-4  | | 3.8e+02| 3.1e+02| 4.6e+02|
NGC1222         |CO6-5  | | 3.1e+02| 2.8e+02| 3.5e+02|
NGC1222         |CO7-6  | | 2.4e+02| 2.2e+02| 2.7e+02|
NGC1222         |CO8-7  | | 1.8e+02| 1.5e+02| 2.2e+02|
NGC1222         |CO9-8  | | 1.0e+02| 4.3e+01| 1.7e+02| 2.6e+02
NGC1222         |CO10-9 | | 6.9e+01| 2.0e+01| 1.1e+02| 2.0e+02
NGC1222         |CO11-10| | 7.3e+01| 3.6e+01| 1.2e+02| 2.0e+02
NGC1222         |CO12-11| | 4.5e+01| 1.3e+01| 8.8e+01| 1.7e+02
NGC1222         |CO13-12| | 9.9e+01| 4.4e+01| 1.5e+02| 2.4e+02
NGC1222         |NII    | | 9.7e+02| 9.2e+02| 1.0e+03|
UGC02608        |CI1-0  | | 3.3e+02| 1.0e+02| 5.0e+02| 7.6e+02
UGC02608        |CI2-1  | | 3.8e+02| 3.2e+02| 4.2e+02|
UGC02608        |CO5-4  | | 1.8e+02| 4.7e+01| 3.1e+02| 5.3e+02
UGC02608        |CO6-5  | | 3.4e+02| 2.7e+02| 4.1e+02|
UGC02608        |CO7-6  | | 1.3e+02| 8.2e+01| 1.8e+02|
UGC02608        |CO9-8  | | 2.1e+02| 8.9e+01| 3.3e+02| 4.7e+02
UGC02608        |CO10-9 | | 1.3e+02| 3.9e+01| 2.1e+02| 3.2e+02
UGC02608        |CO13-12| | 7.8e+01| 2.7e+01| 1.4e+02| 2.3e+02
UGC02608        |NII    | | 1.2e+03| 1.1e+03| 1.3e+03|
NGC1266         |CI1-0  | | 6.8e+02| 4.8e+02| 8.6e+02|
NGC1266         |CI2-1  | | 8.2e+02| 7.7e+02| 8.8e+02|
NGC1266         |CO4-3  | | 1.6e+03| 1.4e+03| 1.8e+03|
NGC1266         |CO5-4  | | 1.4e+03| 1.3e+03| 1.5e+03|
NGC1266         |CO6-5  | | 1.2e+03| 1.2e+03| 1.3e+03|
NGC1266         |CO7-6  | | 1.1e+03| 1.1e+03| 1.2e+03|
NGC1266         |CO8-7  | | 8.8e+02| 8.2e+02| 9.3e+02|
NGC1266         |CO9-8  | | 1.3e+03| 1.2e+03| 1.4e+03|
NGC1266         |CO10-9 | | 9.5e+02| 9.0e+02| 1.0e+03|
NGC1266         |CO11-10| | 9.5e+02| 8.7e+02| 1.0e+03|
NGC1266         |CO12-11| | 6.1e+02| 5.4e+02| 6.7e+02|
NGC1266         |CO13-12| | 2.8e+02| 1.7e+02| 3.8e+02|
NGC1266         |NII    |X| 1.1e+03| 9.5e+02| 1.2e+03|
IRAS 03158+4227 |CI2-1  | | 1.0e+02| 4.3e+01| 1.6e+02|
IRAS 03158+4227 |CO5-4  | | 1.6e+02| 4.0e+01| 3.2e+02| 5.0e+02
IRAS 03158+4227 |CO6-5  | | 2.1e+02| 9.8e+01| 3.3e+02|
IRAS 03158+4227 |CO7-6  | | 2.3e+02| 1.7e+02| 2.9e+02|
IRAS 03158+4227 |CO8-7  | | 1.7e+02| 1.2e+02| 2.2e+02|
IRAS 03158+4227 |CO10-9 | | 1.2e+02| 5.5e+01| 2.1e+02| 3.3e+02
IRAS 03158+4227 |CO11-10| | 1.0e+02| 4.3e+01| 1.5e+02| 2.5e+02
IRAS 03158+4227 |NII    | | 1.0e+02| 3.7e+01| 1.5e+02| 2.3e+02
3C 84           |CI1-0  | | 1.7e+02| 5.8e+01| 2.8e+02| 5.1e+02
3C 84           |CI2-1  | | 4.8e+02| 4.3e+02| 5.1e+02|
3C 84           |CO4-3  | | 3.0e+02| 9.4e+01| 4.4e+02| 7.6e+02
3C 84           |CO5-4  | | 4.7e+02| 3.9e+02| 5.5e+02|
3C 84           |CO6-5  | | 3.7e+02| 3.3e+02| 4.2e+02|
3C 84           |CO7-6  | | 2.7e+02| 2.3e+02| 3.1e+02|
3C 84           |CO8-7  | | 3.0e+02| 2.5e+02| 3.5e+02|
3C 84           |CO9-8  | | 3.4e+02| 2.7e+02| 4.2e+02|
3C 84           |CO10-9 | | 3.6e+02| 3.0e+02| 4.1e+02|
3C 84           |CO11-10| | 2.5e+02| 1.9e+02| 3.0e+02|
3C 84           |CO12-11| | 2.2e+02| 1.7e+02| 2.6e+02|
3C 84           |CO13-12| | 1.3e+02| 7.7e+01| 1.8e+02|
3C 84           |NII    | | 4.6e+02| 4.2e+02| 5.1e+02|
NGC1365-SW      |CI1-0  | | 3.7e+03| 3.4e+03| 4.0e+03|
NGC1365-SW      |CI2-1  | | 4.6e+03| 4.5e+03| 4.8e+03|
NGC1365-SW      |CO4-3  | | 8.0e+03| 7.6e+03| 8.2e+03|
NGC1365-SW      |CO5-4  | | 7.5e+03| 7.4e+03| 7.8e+03|
NGC1365-SW      |CO6-5  | | 5.9e+03| 5.7e+03| 6.0e+03|
NGC1365-SW      |CO7-6  | | 3.7e+03| 3.6e+03| 3.8e+03|
NGC1365-SW      |CO8-7  | | 3.6e+03| 3.2e+03| 3.9e+03|
NGC1365-SW      |CO9-8  | | 1.6e+03| 1.3e+03| 2.0e+03|
NGC1365-SW      |CO10-9 | | 9.8e+02| 7.4e+02| 1.2e+03|
NGC1365-SW      |CO11-10| | 5.1e+02| 2.5e+02| 7.3e+02| 1.1e+03
NGC1365-SW      |CO12-11| | 3.6e+02| 1.5e+02| 5.7e+02| 9.6e+02
NGC1365-SW      |NII    | | 2.1e+04| 2.0e+04| 2.1e+04|
NGC1365-NE      |CI1-0  | | 4.2e+03| 3.8e+03| 4.4e+03|
NGC1365-NE      |CI2-1  | | 4.8e+03| 4.7e+03| 4.9e+03|
NGC1365-NE      |CO4-3  | | 9.1e+03| 8.7e+03| 9.5e+03|
NGC1365-NE      |CO5-4  | | 8.4e+03| 8.1e+03| 8.6e+03|
NGC1365-NE      |CO6-5  | | 6.1e+03| 6.0e+03| 6.2e+03|
NGC1365-NE      |CO7-6  | | 3.8e+03| 3.7e+03| 3.9e+03|
NGC1365-NE      |CO8-7  | | 3.0e+03| 2.7e+03| 3.2e+03|
NGC1365-NE      |CO9-8  | | 1.6e+03| 1.4e+03| 1.8e+03|
NGC1365-NE      |CO10-9 | | 6.3e+02| 4.7e+02| 8.0e+02| 1.1e+03
NGC1365-NE      |CO11-10| | 6.8e+02| 5.6e+02| 8.4e+02|
NGC1365-NE      |CO12-11| | 4.4e+02| 2.5e+02| 5.5e+02| 7.8e+02
NGC1365-NE      |CO13-12| | 2.0e+02| 3.5e+01| 5.0e+02| 9.5e+02
NGC1365-NE      |NII    | | 1.6e+04| 1.6e+04| 1.6e+04|
NGC1377         |CI1-0  | | 2.2e+02| 1.7e+02| 2.8e+02|
NGC1377         |CI2-1  | | 4.5e+01| 2.2e+01| 6.2e+01|
NGC1377         |CO4-3  | | 3.5e+02| 2.7e+02| 4.3e+02|
NGC1377         |CO5-4  | | 1.8e+02| 1.4e+02| 2.4e+02|
NGC1377         |CO6-5  | | 1.3e+02| 1.0e+02| 1.5e+02|
NGC1377         |CO7-6  | | 1.1e+02| 9.0e+01| 1.3e+02|
NGC1377         |CO8-7  | | 2.9e+01| 1.2e+01| 4.7e+01| 8.8e+01
NGC1377         |CO9-8  | | 1.3e+02| 8.5e+01| 1.9e+02|
NGC1377         |CO10-9 | | 1.6e+02| 1.2e+02| 2.0e+02|
NGC1377         |CO11-10| | 1.6e+02| 1.1e+02| 2.1e+02|
NGC1377         |CO12-11| | 1.2e+02| 7.9e+01| 1.6e+02|
NGC1377         |CO13-12| | 2.0e+02| 1.5e+02| 2.4e+02|
NGC1377         |NII    | | 1.5e+02| 1.0e+02| 1.9e+02|
NGC1482         |CI1-0  | | 1.2e+03| 9.6e+02| 1.4e+03|
NGC1482         |CI2-1  | | 1.2e+03| 1.2e+03| 1.3e+03|
NGC1482         |CO4-3  | | 1.7e+03| 1.4e+03| 2.0e+03|
NGC1482         |CO5-4  | | 2.2e+03| 2.0e+03| 2.4e+03|
NGC1482         |CO6-5  | | 1.8e+03| 1.7e+03| 1.9e+03|
NGC1482         |CO7-6  | | 8.7e+02| 8.0e+02| 9.4e+02|
NGC1482         |CO8-7  | | 3.9e+02| 2.6e+02| 5.0e+02|
NGC1482         |CO9-8  | | 4.0e+02| 2.5e+02| 5.4e+02|
NGC1482         |CO10-9 | | 5.5e+02| 4.3e+02| 6.7e+02|
NGC1482         |CO11-10| | 5.1e+02| 3.6e+02| 6.7e+02|
NGC1482         |CO12-11| | 1.5e+02| 5.2e+01| 2.6e+02| 4.2e+02
NGC1482         |CO13-12| | 5.9e+02| 3.2e+02| 8.7e+02|
NGC1482         |NII    | | 6.9e+03| 6.7e+03| 7.2e+03|
IRAS 03521+0028 |CI2-1  | | 3.1e+01| 6.2e+00| 7.8e+01| 1.4e+02
IRAS 03521+0028 |CO5-4  | | 1.5e+02| 4.0e+01| 2.6e+02| 4.6e+02
IRAS 03521+0028 |CO6-5  | | 1.5e+02| 6.5e+01| 2.5e+02| 3.9e+02
IRAS 03521+0028 |CO7-6  | | 8.9e+01| 4.6e+01| 1.5e+02| 2.3e+02
IRAS 03521+0028 |CO8-7  | | 1.3e+02| 8.3e+01| 1.9e+02|
IRAS 03521+0028 |CO10-9 | | 9.9e+01| 6.9e+01| 1.2e+02|
IRAS 03521+0028 |CO11-10| | 3.5e+01| 1.2e+01| 6.8e+01| 9.7e+01
IRAS 03521+0028 |CO12-11| | 2.2e+01| 7.7e+00| 4.3e+01| 6.9e+01
IRAS 03521+0028 |CO13-12| | 3.0e+01| 1.0e+01| 5.0e+01| 8.4e+01
UGC02982        |CI1-0  | | 2.6e+02| 7.0e+01| 4.9e+02| 8.5e+02
UGC02982        |CI2-1  | | 4.3e+02| 3.2e+02| 5.2e+02|
UGC02982        |CO5-4  | | 4.6e+02| 2.6e+02| 6.9e+02| 1.0e+03
UGC02982        |CO6-5  | | 3.8e+02| 2.6e+02| 4.8e+02|
UGC02982        |CO7-6  | | 2.1e+02| 1.0e+02| 3.0e+02| 4.4e+02
UGC02982        |CO8-7  | | 9.7e+01| 2.3e+01| 1.9e+02| 4.4e+02
UGC02982        |CO9-8  | | 1.4e+02| 4.6e+01| 2.6e+02| 4.2e+02
UGC02982        |CO11-10| | 1.3e+02| 4.7e+01| 2.6e+02| 4.4e+02
UGC02982        |CO12-11| | 1.4e+02| 3.6e+01| 2.7e+02| 4.4e+02
UGC02982        |NII    | | 3.1e+03| 3.0e+03| 3.3e+03|
ESO420-G013     |CI1-0  | | 1.2e+03| 5.4e+02| 1.8e+03|
ESO420-G013     |CI2-1  | | 1.0e+03| 8.7e+02| 1.1e+03|
ESO420-G013     |CO4-3  | | 1.9e+03| 1.1e+03| 2.6e+03|
ESO420-G013     |CO5-4  | | 1.5e+03| 1.1e+03| 1.9e+03|
ESO420-G013     |CO6-5  | | 1.2e+03| 9.4e+02| 1.3e+03|
ESO420-G013     |CO7-6  | | 6.6e+02| 5.4e+02| 7.8e+02|
ESO420-G013     |CO8-7  | | 2.7e+02| 8.5e+01| 4.6e+02| 7.7e+02
ESO420-G013     |CO9-8  | | 1.6e+02| 5.0e+01| 3.0e+02| 5.3e+02
ESO420-G013     |CO10-9 | | 1.5e+02| 4.8e+01| 2.8e+02| 5.4e+02
ESO420-G013     |CO11-10| | 9.2e+01| 2.2e+01| 1.8e+02| 3.8e+02
ESO420-G013     |CO12-11| | 3.6e+02| 2.4e+02| 4.7e+02|
ESO420-G013     |CO13-12| | 1.6e+02| 4.3e+01| 3.0e+02| 4.4e+02
ESO420-G013     |NII    | | 2.6e+03| 2.5e+03| 2.8e+03|
NGC1572         |CI1-0  | | 4.8e+02| 1.3e+02| 1.0e+03| 1.7e+03
NGC1572         |CI2-1  | | 9.3e+02| 8.2e+02| 1.0e+03|
NGC1572         |CO5-4  | | 1.4e+03| 1.0e+03| 1.7e+03|
NGC1572         |CO6-5  | | 1.1e+03| 8.7e+02| 1.2e+03|
NGC1572         |CO7-6  | | 7.3e+02| 6.3e+02| 8.4e+02|
NGC1572         |CO8-7  | | 3.6e+02| 2.1e+02| 5.0e+02|
NGC1572         |CO9-8  | | 1.6e+02| 5.1e+01| 2.8e+02| 4.7e+02
NGC1572         |CO10-9 | | 1.2e+02| 3.9e+01| 2.2e+02| 3.8e+02
NGC1572         |CO11-10| | 1.2e+02| 4.0e+01| 2.4e+02| 4.0e+02
NGC1572         |CO12-11| | 1.4e+02| 6.3e+01| 2.4e+02| 3.6e+02
NGC1572         |NII    |X| 2.4e+03| 2.3e+03| 2.6e+03|
IRAS04271+3849  |CI1-0  | | 5.1e+01| 5.5e+00| 1.2e+02| 3.0e+02
IRAS04271+3849  |CI2-1  | | 2.2e+02| 1.8e+02| 2.6e+02|
IRAS04271+3849  |CO5-4  | | 2.5e+02| 1.1e+02| 3.5e+02| 5.2e+02
IRAS04271+3849  |CO6-5  | | 2.5e+02| 2.0e+02| 3.1e+02|
IRAS04271+3849  |CO7-6  | | 1.8e+02| 1.4e+02| 2.2e+02|
IRAS04271+3849  |CO8-7  | | 2.9e+02| 2.1e+02| 3.6e+02|
IRAS04271+3849  |CO9-8  | | 8.6e+01| 2.7e+01| 1.5e+02| 2.7e+02
IRAS04271+3849  |CO10-9 | | 1.7e+02| 9.4e+01| 2.2e+02|
IRAS04271+3849  |CO13-12| | 5.1e+01| 1.4e+01| 9.2e+01| 1.9e+02
IRAS04271+3849  |NII    |X| 1.8e+03| 1.8e+03| 1.9e+03|
NGC1614         |CI1-0  | | 8.4e+02| 5.0e+02| 1.1e+03|
NGC1614         |CI2-1  | | 1.1e+03| 1.0e+03| 1.1e+03|
NGC1614         |CO4-3  | | 2.1e+03| 1.7e+03| 2.4e+03|
NGC1614         |CO5-4  | | 2.2e+03| 2.1e+03| 2.4e+03|
NGC1614         |CO6-5  | | 1.7e+03| 1.6e+03| 1.8e+03|
NGC1614         |CO7-6  | | 1.4e+03| 1.4e+03| 1.5e+03|
NGC1614         |CO8-7  | | 1.1e+03| 1.0e+03| 1.2e+03|
NGC1614         |CO9-8  | | 7.0e+02| 6.3e+02| 7.7e+02|
NGC1614         |CO10-9 | | 5.9e+02| 5.3e+02| 6.6e+02|
NGC1614         |CO11-10| | 2.8e+02| 2.2e+02| 3.4e+02|
NGC1614         |CO12-11| | 2.0e+02| 1.4e+02| 2.5e+02|
NGC1614         |CO13-12| | 1.0e+02| 3.8e+01| 1.7e+02| 2.8e+02
NGC1614         |NII    |X| 2.2e+03| 2.1e+03| 2.3e+03|
UGC03094        |CI1-0  | | 3.2e+02| 1.4e+02| 5.3e+02| 8.3e+02
UGC03094        |CI2-1  | | 3.1e+02| 2.6e+02| 3.6e+02|
UGC03094        |CO5-4  | | 2.1e+02| 8.8e+01| 3.5e+02| 5.4e+02
UGC03094        |CO6-5  | | 2.7e+02| 2.0e+02| 3.4e+02|
UGC03094        |CO7-6  | | 1.1e+02| 6.6e+01| 1.6e+02|
UGC03094        |CO8-7  | | 5.4e+01| 2.0e+01| 1.1e+02| 2.2e+02
UGC03094        |CO9-8  | | 1.2e+02| 4.0e+01| 2.4e+02| 4.6e+02
UGC03094        |CO10-9 | | 2.0e+02| 1.2e+02| 3.1e+02| 4.4e+02
UGC03094        |CO11-10| | 7.8e+01| 2.0e+01| 1.5e+02| 3.0e+02
UGC03094        |NII    | | 1.7e+03| 1.6e+03| 1.8e+03|
MCG-05-12-006   |CI1-0  | | 4.3e+02| 1.5e+02| 7.7e+02| 1.4e+03
MCG-05-12-006   |CI2-1  | | 4.6e+02| 3.6e+02| 5.6e+02|
MCG-05-12-006   |CO5-4  | | 3.9e+02| 1.6e+02| 6.6e+02| 1.1e+03
MCG-05-12-006   |CO6-5  | | 5.0e+02| 3.7e+02| 6.4e+02|
MCG-05-12-006   |CO7-6  | | 6.4e+02| 5.3e+02| 7.3e+02|
MCG-05-12-006   |CO8-7  | | 1.1e+02| 2.9e+01| 2.5e+02| 4.3e+02
MCG-05-12-006   |CO9-8  | | 5.3e+02| 3.3e+02| 7.0e+02|
MCG-05-12-006   |CO10-9 | | 3.3e+02| 2.3e+02| 4.7e+02|
MCG-05-12-006   |CO12-11| | 8.3e+01| 1.6e+01| 1.6e+02| 3.4e+02
MCG-05-12-006   |NII    | | 7.2e+02| 6.2e+02| 8.2e+02|
IRAS F05189-2524|CI1-0  | | 3.6e+02| 1.5e+02| 5.6e+02| 7.7e+02
IRAS F05189-2524|CI2-1  | | 2.1e+02| 1.6e+02| 2.6e+02|
IRAS F05189-2524|CO5-4  | | 2.6e+02| 1.2e+02| 3.8e+02| 6.0e+02
IRAS F05189-2524|CO6-5  | | 3.8e+02| 3.1e+02| 4.5e+02|
IRAS F05189-2524|CO7-6  | | 3.0e+02| 2.4e+02| 3.5e+02|
IRAS F05189-2524|CO8-7  | | 3.9e+02| 3.3e+02| 4.4e+02|
IRAS F05189-2524|CO9-8  | | 2.3e+02| 1.8e+02| 2.7e+02|
IRAS F05189-2524|CO10-9 | | 2.6e+02| 2.2e+02| 2.9e+02|
IRAS F05189-2524|CO11-10| | 1.6e+02| 1.3e+02| 1.9e+02|
IRAS F05189-2524|CO12-11| | 1.5e+02| 1.2e+02| 1.7e+02|
IRAS F05189-2524|CO13-12| | 1.4e+02| 1.1e+02| 1.6e+02|
IRAS F05189-2524|NII    | | 1.9e+02| 1.6e+02| 2.1e+02|
IRAS05223+1908  |CO7-6  | | 1.7e+02| 1.7e+02| 1.7e+02|
IRAS05223+1908  |CO8-7  | | 8.1e+01| 8.1e+01| 8.1e+01|
MCG+08-11-002   |CI1-0  | | 8.2e+02| 4.3e+02| 1.3e+03|
MCG+08-11-002   |CI2-1  | | 1.0e+03| 9.3e+02| 1.1e+03|
MCG+08-11-002   |CO5-4  | | 1.6e+03| 1.4e+03| 2.0e+03|
MCG+08-11-002   |CO6-5  | | 1.2e+03| 1.1e+03| 1.3e+03|
MCG+08-11-002   |CO7-6  | | 8.0e+02| 7.0e+02| 8.8e+02|
MCG+08-11-002   |CO8-7  | | 6.0e+02| 4.8e+02| 7.2e+02|
MCG+08-11-002   |CO9-8  | | 5.6e+02| 4.3e+02| 7.0e+02|
MCG+08-11-002   |CO10-9 | | 3.0e+02| 2.1e+02| 4.1e+02|
MCG+08-11-002   |CO11-10| | 1.9e+02| 8.2e+01| 2.8e+02| 4.4e+02
MCG+08-11-002   |CO12-11| | 7.9e+01| 2.3e+01| 1.5e+02| 2.6e+02
MCG+08-11-002   |CO13-12| | 1.5e+02| 5.2e+01| 2.3e+02| 3.8e+02
MCG+08-11-002   |NII    | | 1.1e+03| 1.0e+03| 1.2e+03|
NGC1961         |CI1-0  | | 5.0e+02| 2.8e+02| 8.7e+02|
NGC1961         |CI2-1  | | 7.3e+02| 6.3e+02| 8.2e+02|
NGC1961         |CO4-3  | | 1.5e+03| 1.2e+03| 2.0e+03|
NGC1961         |CO5-4  | | 1.1e+03| 9.2e+02| 1.3e+03|
NGC1961         |CO6-5  | | 5.4e+02| 4.2e+02| 6.6e+02|
NGC1961         |CO7-6  | | 4.9e+02| 3.9e+02| 5.9e+02|
NGC1961         |CO8-7  | | 5.2e+02| 3.7e+02| 6.8e+02|
NGC1961         |CO9-8  | | 3.9e+02| 1.4e+02| 6.7e+02| 1.0e+03
NGC1961         |CO10-9 | | 2.0e+02| 4.4e+01| 4.8e+02| 6.9e+02
NGC1961         |CO11-10| | 2.2e+02| 5.8e+01| 4.4e+02| 7.7e+02
NGC1961         |CO12-11| | 5.0e+02| 3.1e+02| 7.3e+02|
NGC1961         |CO13-12| | 2.2e+02| 7.2e+01| 4.3e+02| 7.6e+02
NGC1961         |NII    |X| 3.3e+03| 2.8e+03| 3.7e+03|
UGC03351        |CI1-0  | | 6.1e+02| 2.6e+02| 9.6e+02| 1.5e+03
UGC03351        |CI2-1  | | 8.6e+02| 7.6e+02| 9.7e+02|
UGC03351        |CO4-3  | | 1.4e+03| 8.5e+02| 1.9e+03|
UGC03351        |CO5-4  | | 1.2e+03| 8.8e+02| 1.5e+03|
UGC03351        |CO6-5  | | 9.5e+02| 8.1e+02| 1.0e+03|
UGC03351        |CO7-6  | | 5.1e+02| 4.1e+02| 6.2e+02|
UGC03351        |CO8-7  | | 2.6e+02| 1.1e+02| 3.8e+02| 5.8e+02
UGC03351        |CO9-8  | | 1.4e+02| 4.0e+01| 2.7e+02| 5.1e+02
UGC03351        |CO10-9 | | 2.6e+02| 1.3e+02| 4.0e+02| 6.0e+02
UGC03351        |CO11-10| | 1.4e+02| 3.9e+01| 2.7e+02| 4.5e+02
UGC03351        |CO13-12| | 1.8e+02| 8.8e+01| 2.9e+02| 4.8e+02
UGC03351        |NII    | | 2.2e+03| 2.1e+03| 2.3e+03|
IRAS05442+1732  |CI1-0  | | 6.4e+02| 2.7e+02| 1.2e+03| 2.0e+03
IRAS05442+1732  |CI2-1  | | 3.3e+02| 2.4e+02| 4.1e+02|
IRAS05442+1732  |CO5-4  | | 6.6e+02| 2.8e+02| 1.1e+03| 1.8e+03
IRAS05442+1732  |CO6-5  | | 5.1e+02| 3.9e+02| 6.9e+02|
IRAS05442+1732  |CO7-6  | | 3.8e+02| 2.9e+02| 4.6e+02|
IRAS05442+1732  |CO8-7  | | 4.5e+02| 3.4e+02| 5.4e+02|
IRAS05442+1732  |CO9-8  | | 2.4e+02| 1.0e+02| 3.9e+02| 6.0e+02
IRAS05442+1732  |CO11-10| | 1.6e+02| 4.0e+01| 2.6e+02| 4.6e+02
IRAS05442+1732  |CO13-12| | 1.2e+02| 4.7e+01| 2.2e+02| 3.4e+02
IRAS05442+1732  |NII    | | 7.1e+02| 6.3e+02| 7.9e+02|
IRAS 06035-7102 |CI1-0  | | 1.1e+02| 1.1e+01| 2.4e+02| 4.4e+02
IRAS 06035-7102 |CI2-1  | | 1.5e+02| 1.0e+02| 2.0e+02|
IRAS 06035-7102 |CO5-4  | | 5.2e+02| 3.2e+02| 6.8e+02|
IRAS 06035-7102 |CO6-5  | | 2.7e+02| 1.8e+02| 3.6e+02|
IRAS 06035-7102 |CO7-6  | | 3.1e+02| 2.6e+02| 3.6e+02|
IRAS 06035-7102 |CO8-7  | | 3.3e+02| 2.8e+02| 3.8e+02|
IRAS 06035-7102 |CO9-8  | | 2.8e+02| 2.2e+02| 3.6e+02|
IRAS 06035-7102 |CO10-9 | | 3.0e+02| 2.5e+02| 3.6e+02|
IRAS 06035-7102 |CO11-10| | 2.2e+02| 1.8e+02| 2.6e+02|
IRAS 06035-7102 |CO12-11| | 1.4e+02| 9.1e+01| 1.9e+02|
IRAS 06035-7102 |CO13-12| | 3.6e+01| 1.0e+01| 7.1e+01| 1.3e+02
IRAS 06035-7102 |NII    | | 2.5e+02| 2.1e+02| 2.9e+02|
UGC03410a       |CI1-0  | | 5.9e+02| 2.3e+02| 9.0e+02| 1.3e+03
UGC03410a       |CI2-1  | | 5.8e+02| 4.8e+02| 6.8e+02|
UGC03410a       |CO4-3  | | 4.2e+02| 1.1e+02| 8.5e+02| 1.6e+03
UGC03410a       |CO5-4  | | 3.3e+02| 1.3e+02| 5.3e+02| 8.8e+02
UGC03410a       |CO6-5  | | 3.4e+02| 2.3e+02| 4.6e+02|
UGC03410a       |CO7-6  | | 6.6e+01| 1.2e+01| 1.5e+02| 2.4e+02
UGC03410a       |CO9-8  | | 2.3e+02| 7.6e+01| 4.1e+02| 7.6e+02
UGC03410a       |CO10-9 | | 1.3e+02| 2.5e+01| 2.8e+02| 5.2e+02
UGC03410a       |CO11-10| | 3.0e+02| 1.1e+02| 4.5e+02| 7.2e+02
UGC03410a       |CO13-12| | 2.1e+02| 6.4e+01| 3.8e+02| 6.4e+02
UGC03410a       |NII    | | 4.1e+03| 3.9e+03| 4.3e+03|
NGC2146-NW      |CI1-0  | | 3.3e+03| 3.0e+03| 3.5e+03|
NGC2146-NW      |CI2-1  | | 4.1e+03| 4.0e+03| 4.2e+03|
NGC2146-NW      |CO4-3  | | 7.6e+03| 7.2e+03| 8.0e+03|
NGC2146-NW      |CO5-4  | | 7.4e+03| 7.2e+03| 7.6e+03|
NGC2146-NW      |CO6-5  | | 6.7e+03| 6.6e+03| 6.8e+03|
NGC2146-NW      |CO7-6  | | 4.5e+03| 4.3e+03| 4.6e+03|
NGC2146-NW      |CO8-7  | | 3.4e+03| 3.2e+03| 3.6e+03|
NGC2146-NW      |CO9-8  | | 2.3e+03| 2.0e+03| 2.6e+03|
NGC2146-NW      |CO10-9 | | 9.8e+02| 7.9e+02| 1.2e+03|
NGC2146-NW      |CO11-10| | 7.0e+02| 5.0e+02| 9.2e+02|
NGC2146-NW      |CO12-11| | 6.4e+02| 4.5e+02| 8.1e+02|
NGC2146-NW      |NII    | | 1.9e+04| 1.9e+04| 2.0e+04|
NGC2146-nuc     |CI1-0  | | 2.6e+03| 2.3e+03| 2.9e+03|
NGC2146-nuc     |CI2-1  | | 4.6e+03| 4.5e+03| 4.7e+03|
NGC2146-nuc     |CO4-3  | | 7.7e+03| 7.3e+03| 8.1e+03|
NGC2146-nuc     |CO5-4  | | 8.3e+03| 8.1e+03| 8.5e+03|
NGC2146-nuc     |CO6-5  | | 7.5e+03| 7.4e+03| 7.6e+03|
NGC2146-nuc     |CO7-6  | | 5.4e+03| 5.3e+03| 5.5e+03|
NGC2146-nuc     |CO8-7  | | 4.4e+03| 4.2e+03| 4.5e+03|
NGC2146-nuc     |CO9-8  | | 2.9e+03| 2.7e+03| 3.1e+03|
NGC2146-nuc     |CO10-9 | | 1.8e+03| 1.6e+03| 2.0e+03|
NGC2146-nuc     |CO11-10| | 1.2e+03| 1.0e+03| 1.5e+03|
NGC2146-nuc     |CO12-11| | 5.2e+02| 3.2e+02| 7.2e+02| 9.6e+02
NGC2146-nuc     |CO13-12| | 5.6e+02| 2.2e+02| 9.6e+02| 1.5e+03
NGC2146-nuc     |NII    | | 2.7e+04| 2.6e+04| 2.7e+04|
NGC2146-SE      |CI1-0  | | 2.8e+03| 2.5e+03| 3.2e+03|
NGC2146-SE      |CI2-1  | | 3.9e+03| 3.8e+03| 4.0e+03|
NGC2146-SE      |CO4-3  | | 7.4e+03| 7.0e+03| 7.8e+03|
NGC2146-SE      |CO5-4  | | 7.0e+03| 6.7e+03| 7.2e+03|
NGC2146-SE      |CO6-5  | | 6.6e+03| 6.5e+03| 6.8e+03|
NGC2146-SE      |CO7-6  | | 4.7e+03| 4.6e+03| 4.8e+03|
NGC2146-SE      |CO8-7  | | 3.8e+03| 3.6e+03| 4.0e+03|
NGC2146-SE      |CO9-8  | | 2.2e+03| 1.9e+03| 2.5e+03|
NGC2146-SE      |CO10-9 | | 1.3e+03| 1.0e+03| 1.5e+03|
NGC2146-SE      |CO11-10| | 1.0e+03| 7.5e+02| 1.2e+03|
NGC2146-SE      |CO12-11| | 4.0e+02| 1.6e+02| 6.4e+02| 1.0e+03
NGC2146-SE      |CO13-12| | 6.6e+02| 2.3e+02| 1.2e+03| 2.0e+03
NGC2146-SE      |NII    | | 2.2e+04| 2.1e+04| 2.2e+04|
IRAS 06206-6315 |CI2-1  | | 1.4e+02| 9.9e+01| 1.9e+02|
IRAS 06206-6315 |CO5-4  | | 1.7e+02| 4.6e+01| 2.8e+02| 4.0e+02
IRAS 06206-6315 |CO6-5  | | 1.8e+02| 9.7e+01| 2.7e+02| 3.7e+02
IRAS 06206-6315 |CO7-6  | | 1.8e+02| 1.3e+02| 2.2e+02|
IRAS 06206-6315 |CO8-7  | | 1.4e+02| 1.0e+02| 1.8e+02|
IRAS 06206-6315 |CO10-9 | | 8.3e+01| 4.3e+01| 1.2e+02| 1.8e+02
IRAS 06206-6315 |CO11-10| | 7.9e+01| 4.2e+01| 1.2e+02| 1.7e+02
IRAS 06206-6315 |CO12-11| | 2.9e+01| 6.5e+00| 5.4e+01| 8.8e+01
IRAS 06206-6315 |NII    | | 8.0e+01| 4.8e+01| 1.1e+02|
ESO255-IG007    |CI1-0  | | 3.4e+02| 1.2e+02| 6.3e+02| 1.0e+03
ESO255-IG007    |CI2-1  | | 3.7e+02| 3.2e+02| 4.2e+02|
ESO255-IG007    |CO5-4  | | 5.1e+02| 3.0e+02| 6.7e+02| 8.9e+02
ESO255-IG007    |CO6-5  | | 4.7e+02| 3.7e+02| 5.5e+02|
ESO255-IG007    |CO7-6  | | 3.2e+02| 2.6e+02| 3.8e+02|
ESO255-IG007    |CO8-7  | | 3.0e+02| 2.3e+02| 3.7e+02|
ESO255-IG007    |CO9-8  | | 2.9e+02| 2.2e+02| 3.5e+02|
ESO255-IG007    |CO10-9 | | 2.2e+02| 1.6e+02| 2.6e+02|
ESO255-IG007    |CO12-11| | 4.0e+01| 7.0e+00| 7.8e+01| 1.5e+02
ESO255-IG007    |CO13-12| | 7.0e+01| 2.8e+01| 1.2e+02| 1.8e+02
ESO255-IG007    |NII    | | 6.1e+02| 5.6e+02| 6.6e+02|
UGC03608        |CI1-0  | | 2.9e+02| 9.9e+01| 4.7e+02| 7.8e+02
UGC03608        |CI2-1  | | 4.5e+02| 3.9e+02| 5.0e+02|
UGC03608        |CO5-4  | | 8.6e+02| 7.0e+02| 9.9e+02|
UGC03608        |CO6-5  | | 4.9e+02| 4.4e+02| 5.6e+02|
UGC03608        |CO7-6  | | 3.8e+02| 3.3e+02| 4.4e+02|
UGC03608        |CO8-7  | | 3.0e+02| 2.3e+02| 3.7e+02|
UGC03608        |CO9-8  | | 2.0e+02| 6.1e+01| 3.1e+02| 5.1e+02
UGC03608        |CO10-9 | | 1.7e+02| 7.1e+01| 2.6e+02| 4.1e+02
UGC03608        |CO11-10| | 8.6e+01| 1.5e+01| 1.9e+02| 2.8e+02
UGC03608        |CO12-11| | 9.2e+01| 3.3e+01| 1.6e+02| 2.7e+02
UGC03608        |CO13-12| | 2.9e+01| 2.0e+00| 9.6e+01| 2.2e+02
UGC03608        |NII    | | 1.2e+03| 1.1e+03| 1.2e+03|
NGC2342b        |CI1-0  | | 1.9e+02| 4.0e+01| 3.6e+02| 8.7e+02
NGC2342b        |CI2-1  | | 3.4e+02| 2.8e+02| 4.0e+02|
NGC2342b        |CO4-3  | | 4.7e+02| 1.6e+02| 8.6e+02| 1.7e+03
NGC2342b        |CO5-4  | | 3.8e+02| 1.4e+02| 5.6e+02| 8.5e+02
NGC2342b        |CO6-5  | | 2.9e+02| 1.8e+02| 4.0e+02|
NGC2342b        |CO7-6  | | 2.6e+02| 2.1e+02| 3.2e+02|
NGC2342b        |CO8-7  | | 2.8e+02| 1.8e+02| 3.4e+02|
NGC2342b        |CO10-9 | | 9.4e+01| 2.3e+01| 1.7e+02| 3.0e+02
NGC2342b        |CO12-11| | 1.6e+02| 8.9e+01| 2.3e+02| 3.4e+02
NGC2342b        |CO13-12| | 7.3e+01| 1.5e+01| 1.4e+02| 2.5e+02
NGC2342b        |NII    | | 1.7e+03| 1.6e+03| 1.8e+03|
NGC2342a        |CI1-0  | | 5.6e+02| 2.8e+02| 8.1e+02| 1.2e+03
NGC2342a        |CI2-1  | | 3.8e+02| 3.2e+02| 4.4e+02|
NGC2342a        |CO4-3  | | 1.0e+03| 7.5e+02| 1.3e+03|
NGC2342a        |CO6-5  | | 4.8e+02| 3.8e+02| 5.8e+02|
NGC2342a        |CO7-6  | | 2.4e+02| 1.8e+02| 3.0e+02|
NGC2342a        |CO8-7  | | 1.6e+02| 5.8e+01| 2.5e+02| 4.4e+02
NGC2342a        |CO9-8  | | 6.2e+01| 6.8e+00| 1.8e+02| 4.2e+02
NGC2342a        |CO10-9 | | 1.8e+02| 3.9e+01| 3.2e+02| 5.1e+02
NGC2342a        |CO13-12| | 2.1e+02| 6.6e+01| 3.6e+02| 5.8e+02
NGC2342a        |NII    | | 1.4e+03| 1.3e+03| 1.6e+03|
NGC2369         |CI1-0  | | 1.4e+03| 8.7e+02| 1.8e+03|
NGC2369         |CI2-1  | | 1.4e+03| 1.3e+03| 1.6e+03|
NGC2369         |CO4-3  | | 1.4e+03| 7.2e+02| 1.8e+03| 2.6e+03
NGC2369         |CO5-4  | | 2.3e+03| 2.0e+03| 2.5e+03|
NGC2369         |CO6-5  | | 1.8e+03| 1.7e+03| 2.0e+03|
NGC2369         |CO7-6  | | 1.2e+03| 1.1e+03| 1.3e+03|
NGC2369         |CO8-7  | | 9.5e+02| 8.2e+02| 1.1e+03|
NGC2369         |CO9-8  | | 6.7e+02| 5.2e+02| 8.6e+02|
NGC2369         |CO10-9 | | 4.2e+02| 2.8e+02| 5.6e+02|
NGC2369         |CO11-10| | 2.6e+02| 1.4e+02| 4.0e+02| 6.3e+02
NGC2369         |CO12-11| | 2.9e+02| 1.9e+02| 4.2e+02|
NGC2369         |CO13-12| | 1.2e+02| 2.7e+01| 2.4e+02| 3.6e+02
NGC2369         |NII    |X| 5.8e+03| 5.7e+03| 6.0e+03|
NGC2388a        |CI1-0  | | 3.2e+02| 1.3e+02| 7.0e+02| 1.2e+03
NGC2388a        |CI2-1  | | 6.9e+02| 6.1e+02| 7.6e+02|
NGC2388a        |CO4-3  | | 7.8e+02| 4.0e+02| 1.2e+03| 1.9e+03
NGC2388a        |CO5-4  | | 7.4e+02| 5.2e+02| 9.7e+02|
NGC2388a        |CO6-5  | | 1.0e+03| 9.1e+02| 1.1e+03|
NGC2388a        |CO7-6  | | 6.9e+02| 6.1e+02| 7.6e+02|
NGC2388a        |CO8-7  | | 5.8e+02| 4.6e+02| 7.0e+02|
NGC2388a        |CO9-8  | | 3.2e+02| 2.2e+02| 4.8e+02|
NGC2388a        |CO10-9 | | 1.2e+02| 2.6e+01| 2.1e+02| 3.2e+02
NGC2388a        |CO11-10| | 9.3e+01| 1.6e+01| 1.8e+02| 3.6e+02
NGC2388a        |CO12-11| | 5.2e+01| 9.4e+00| 1.3e+02| 2.2e+02
NGC2388a        |CO13-12| | 2.3e+02| 1.2e+02| 3.3e+02| 4.8e+02
NGC2388a        |NII    | | 2.1e+03| 2.0e+03| 2.2e+03|
MCG+02-20-003   |CI1-0  | | 3.1e+02| 1.1e+02| 6.1e+02| 1.0e+03
MCG+02-20-003   |CI2-1  | | 3.2e+02| 2.6e+02| 4.0e+02|
MCG+02-20-003   |CO4-3  | | 3.5e+02| 1.1e+02| 7.5e+02| 1.5e+03
MCG+02-20-003   |CO5-4  | | 5.9e+02| 3.6e+02| 7.9e+02|
MCG+02-20-003   |CO6-5  | | 5.4e+02| 4.3e+02| 6.3e+02|
MCG+02-20-003   |CO7-6  | | 2.6e+02| 2.1e+02| 3.4e+02|
MCG+02-20-003   |CO8-7  | | 2.2e+02| 1.3e+02| 3.0e+02| 4.2e+02
MCG+02-20-003   |CO9-8  | | 2.4e+02| 1.4e+02| 3.4e+02|
MCG+02-20-003   |CO10-9 | | 8.0e+01| 3.1e+01| 1.4e+02| 2.6e+02
MCG+02-20-003   |CO11-10| | 2.4e+02| 1.5e+02| 3.1e+02|
MCG+02-20-003   |CO12-11| | 9.8e+01| 3.8e+01| 1.6e+02| 2.5e+02
MCG+02-20-003   |CO13-12| | 6.7e+01| 1.7e+01| 1.2e+02| 1.9e+02
MCG+02-20-003   |NII    | | 7.4e+02| 6.7e+02| 8.0e+02|
IRAS 07598+6508 |CI2-1  | | 3.9e+01| 1.4e+01| 7.0e+01| 1.3e+02
IRAS 07598+6508 |CO5-4  | | 1.1e+02| 3.0e+01| 2.5e+02| 4.2e+02
IRAS 07598+6508 |CO6-5  | | 1.3e+02| 4.9e+01| 2.2e+02| 3.4e+02
IRAS 07598+6508 |CO7-6  | | 4.3e+01| 1.6e+01| 8.4e+01| 1.4e+02
IRAS 07598+6508 |CO8-7  | | 2.9e+01| 8.6e+00| 5.5e+01| 9.0e+01
IRAS 07598+6508 |CO10-9 | | 7.2e+01| 2.0e+01| 1.3e+02| 2.0e+02
IRAS 07598+6508 |CO11-10| | 6.3e+01| 2.1e+01| 1.1e+02| 1.6e+02
IRAS 07598+6508 |CO12-11| | 6.8e+01| 3.3e+01| 1.1e+02| 1.6e+02
IRAS 07598+6508 |CO13-12| | 4.3e+01| 8.8e+00| 7.8e+01| 1.4e+02
IRAS 07598+6508 |NII    | | 5.8e+01| 2.2e+01| 9.5e+01| 1.5e+02
B2 0827+24      |CO8-7  | | 7.9e+01| 2.0e+01| 1.6e+02| 3.5e+02
IRAS 08311-2459 |CI2-1  | | 1.9e+02| 1.4e+02| 2.4e+02|
IRAS 08311-2459 |CO5-4  | | 5.6e+02| 3.4e+02| 7.5e+02|
IRAS 08311-2459 |CO6-5  | | 5.7e+02| 4.8e+02| 6.7e+02|
IRAS 08311-2459 |CO7-6  | | 3.6e+02| 3.2e+02| 4.1e+02|
IRAS 08311-2459 |CO8-7  | | 3.0e+02| 2.5e+02| 3.6e+02|
IRAS 08311-2459 |CO10-9 | | 1.8e+02| 1.4e+02| 2.3e+02|
IRAS 08311-2459 |CO11-10| | 1.4e+02| 8.9e+01| 1.8e+02|
IRAS 08311-2459 |CO12-11| | 1.7e+02| 1.2e+02| 2.0e+02|
IRAS 08311-2459 |CO13-12| | 3.6e+01| 1.0e+01| 6.7e+01| 1.2e+02
IRAS 08311-2459 |NII    | | 2.1e+02| 1.7e+02| 2.4e+02|
He2-10          |CI1-0  | | 2.3e+02| 8.3e+01| 4.1e+02| 5.6e+02
He2-10          |CI2-1  | | 3.1e+02| 2.5e+02| 3.5e+02|
He2-10          |CO4-3  | | 3.6e+02| 2.0e+02| 5.5e+02|
He2-10          |CO5-4  | | 5.5e+02| 4.4e+02| 6.7e+02|
He2-10          |CO6-5  | | 6.0e+02| 5.5e+02| 6.6e+02|
He2-10          |CO7-6  | | 4.6e+02| 4.0e+02| 5.0e+02|
He2-10          |CO8-7  | | 3.5e+02| 2.9e+02| 4.2e+02|
He2-10          |CO9-8  | | 4.0e+02| 3.1e+02| 5.0e+02|
He2-10          |CO10-9 | | 2.6e+02| 1.6e+02| 3.5e+02| 4.8e+02
He2-10          |CO11-10| | 1.4e+02| 6.8e+01| 2.4e+02| 3.4e+02
He2-10          |CO13-12| | 2.4e+02| 1.0e+02| 3.7e+02|
He2-10          |NII    | | 2.1e+03| 2.0e+03| 2.2e+03|
IRAS08355-4944  |CI1-0  | | 8.3e+01| 1.8e+01| 1.6e+02| 2.8e+02
IRAS08355-4944  |CI2-1  | | 9.2e+01| 6.5e+01| 1.2e+02|
IRAS08355-4944  |CO5-4  | | 4.2e+01| 5.1e+00| 9.7e+01| 1.6e+02
IRAS08355-4944  |CO6-5  | | 9.4e+01| 5.3e+01| 1.2e+02| 1.7e+02
IRAS08355-4944  |CO7-6  | | 1.7e+02| 1.5e+02| 1.9e+02|
IRAS08355-4944  |CO8-7  | | 1.9e+02| 1.5e+02| 2.3e+02|
IRAS08355-4944  |CO9-8  | | 1.6e+02| 9.7e+01| 2.4e+02| 3.7e+02
IRAS08355-4944  |CO10-9 | | 3.1e+02| 2.6e+02| 3.6e+02|
IRAS08355-4944  |CO11-10| | 1.3e+02| 6.9e+01| 1.9e+02| 2.8e+02
IRAS08355-4944  |CO12-11| | 1.3e+02| 8.6e+01| 1.9e+02|
IRAS08355-4944  |CO13-12| | 3.6e+02| 2.9e+02| 4.0e+02|
IRAS08355-4944  |NII    | | 5.0e+02| 4.4e+02| 5.5e+02|
NGC2623         |CI1-0  | | 5.4e+02| 3.2e+02| 7.4e+02|
NGC2623         |CI2-1  | | 7.5e+02| 7.0e+02| 7.9e+02|
NGC2623         |CO5-4  | | 1.0e+03| 9.1e+02| 1.1e+03|
NGC2623         |CO6-5  | | 9.6e+02| 9.1e+02| 1.0e+03|
NGC2623         |CO7-6  | | 8.8e+02| 8.3e+02| 9.2e+02|
NGC2623         |CO8-7  | | 8.8e+02| 8.3e+02| 9.4e+02|
NGC2623         |CO9-8  | | 6.9e+02| 6.4e+02| 7.5e+02|
NGC2623         |CO10-9 | | 6.8e+02| 6.2e+02| 7.4e+02|
NGC2623         |CO11-10| | 4.5e+02| 4.1e+02| 5.0e+02|
NGC2623         |CO12-11| | 3.2e+02| 2.9e+02| 3.5e+02|
NGC2623         |CO13-12| | 2.7e+02| 2.2e+02| 3.1e+02|
NGC2623         |NII    | | 4.4e+02| 3.9e+02| 4.8e+02|
IRAS 08572+3915 |CI1-0  | | 4.1e+02| 1.7e+02| 6.7e+02| 1.1e+03
IRAS 08572+3915 |CI2-1  | | 4.7e+01| 1.4e+01| 8.8e+01| 1.8e+02
IRAS 08572+3915 |CO5-4  | | 1.7e+02| 5.0e+01| 3.0e+02| 5.2e+02
IRAS 08572+3915 |CO6-5  | | 1.5e+02| 7.5e+01| 2.2e+02| 3.6e+02
IRAS 08572+3915 |CO8-7  | | 1.0e+02| 4.8e+01| 1.6e+02| 2.3e+02
IRAS 08572+3915 |CO9-8  | | 8.4e+01| 2.6e+01| 1.7e+02| 3.4e+02
IRAS 08572+3915 |CO10-9 | | 1.2e+02| 5.9e+01| 1.8e+02|
IRAS 08572+3915 |CO11-10| | 1.3e+02| 8.2e+01| 2.0e+02|
IRAS 08572+3915 |CO12-11| | 6.1e+01| 1.8e+01| 1.3e+02| 2.0e+02
IRAS 08572+3915 |CO13-12| | 4.1e+01| 8.8e+00| 7.2e+01| 1.2e+02
IRAS09022-3615  |CI1-0  | | 6.3e+02| 3.7e+02| 8.5e+02| 1.1e+03
IRAS09022-3615  |CI2-1  | | 3.8e+02| 3.4e+02| 4.1e+02|
IRAS09022-3615  |CO5-4  | | 8.0e+02| 6.3e+02| 9.5e+02|
IRAS09022-3615  |CO6-5  | | 6.9e+02| 6.4e+02| 7.6e+02|
IRAS09022-3615  |CO7-6  | | 5.4e+02| 5.1e+02| 5.7e+02|
IRAS09022-3615  |CO8-7  | | 3.4e+02| 3.1e+02| 3.7e+02|
IRAS09022-3615  |CO9-8  | | 4.0e+02| 3.4e+02| 4.6e+02|
IRAS09022-3615  |CO10-9 | | 2.7e+02| 2.4e+02| 3.1e+02|
IRAS09022-3615  |CO11-10| | 2.3e+02| 1.9e+02| 2.7e+02|
IRAS09022-3615  |CO12-11| | 1.6e+02| 1.3e+02| 2.0e+02|
IRAS09022-3615  |CO13-12| | 1.1e+02| 8.4e+01| 1.5e+02|
IRAS09022-3615  |NII    |X| 6.1e+02| 5.6e+02| 6.6e+02|
NGC2764         |CI1-0  | | 4.2e+02| 1.8e+02| 6.4e+02| 9.8e+02
NGC2764         |CI2-1  | | 2.3e+02| 1.9e+02| 2.8e+02|
NGC2764         |CO4-3  | | 1.5e+03| 1.2e+03| 1.8e+03|
NGC2764         |CO5-4  | | 5.3e+02| 3.4e+02| 6.9e+02| 8.9e+02
NGC2764         |CO6-5  | | 1.8e+02| 1.2e+02| 2.5e+02|
NGC2764         |CO7-6  | | 1.4e+02| 9.2e+01| 1.8e+02|
NGC2764         |CO8-7  | | 8.8e+01| 3.7e+01| 1.3e+02| 1.9e+02
NGC2764         |CO9-8  | | 7.4e+01| 1.9e+01| 1.5e+02| 2.6e+02
NGC2764         |CO10-9 | | 6.9e+01| 2.1e+01| 1.3e+02| 2.0e+02
NGC2764         |CO11-10| | 8.5e+01| 3.2e+01| 1.5e+02| 2.6e+02
NGC2764         |CO13-12| | 5.4e+01| 1.3e+01| 1.1e+02| 1.7e+02
NGC2764         |NII    | | 1.4e+03| 1.3e+03| 1.4e+03|
NGC2798         |CI1-0  | | 8.5e+02| 6.8e+02| 1.1e+03|
NGC2798         |CI2-1  | | 8.2e+02| 7.4e+02| 8.8e+02|
NGC2798         |CO4-3  | | 1.7e+03| 1.5e+03| 2.0e+03|
NGC2798         |CO5-4  | | 1.5e+03| 1.4e+03| 1.6e+03|
NGC2798         |CO6-5  | | 1.4e+03| 1.4e+03| 1.5e+03|
NGC2798         |CO7-6  | | 1.1e+03| 9.9e+02| 1.1e+03|
NGC2798         |CO8-7  | | 6.7e+02| 5.8e+02| 7.5e+02|
NGC2798         |CO9-8  | | 5.8e+02| 4.7e+02| 6.8e+02|
NGC2798         |CO10-9 | | 5.2e+02| 4.2e+02| 6.2e+02|
NGC2798         |CO11-10| | 3.8e+02| 3.1e+02| 4.8e+02|
NGC2798         |CO12-11| | 1.5e+02| 7.9e+01| 2.2e+02| 3.2e+02
NGC2798         |CO13-12| | 4.5e+02| 3.0e+02| 5.7e+02|
NGC2798         |NII    |X| 3.7e+03| 3.6e+03| 3.9e+03|
UGC05101        |CI1-0  | | 3.8e+02| 1.6e+02| 6.5e+02| 1.0e+03
UGC05101        |CI2-1  | | 5.1e+02| 4.5e+02| 5.7e+02|
UGC05101        |CO5-4  | | 5.6e+02| 3.7e+02| 7.3e+02|
UGC05101        |CO6-5  | | 5.9e+02| 4.9e+02| 6.8e+02|
UGC05101        |CO7-6  | | 3.7e+02| 3.1e+02| 4.4e+02|
UGC05101        |CO8-7  | | 3.6e+02| 3.0e+02| 4.2e+02|
UGC05101        |CO9-8  | | 2.4e+02| 1.4e+02| 3.4e+02|
UGC05101        |CO10-9 | | 3.1e+02| 2.4e+02| 3.7e+02|
UGC05101        |CO11-10| | 1.7e+02| 9.7e+01| 2.4e+02|
UGC05101        |CO12-11| | 6.5e+01| 1.7e+01| 1.2e+02| 2.0e+02
UGC05101        |CO13-12| | 8.8e+01| 2.8e+01| 1.6e+02| 2.2e+02
UGC05101        |NII    |X| 1.2e+03| 1.2e+03| 1.3e+03|
NGC2976_00      |CI1-0  | | 1.4e+02| 5.3e+01| 2.6e+02| 4.0e+02
NGC2976_00      |CI2-1  | | 6.2e+01| 1.9e+01| 1.1e+02| 2.0e+02
NGC2976_00      |CO4-3  | | 2.5e+02| 5.2e+01| 3.8e+02| 6.4e+02
NGC2976_00      |CO5-4  | | 1.6e+02| 3.8e+01| 3.1e+02| 4.4e+02
NGC2976_00      |CO6-5  | | 8.0e+01| 2.8e+01| 1.6e+02| 2.3e+02
NGC2976_00      |CO7-6  | | 1.2e+02| 6.7e+01| 1.6e+02| 2.2e+02
NGC2976_00      |CO9-8  | | 1.6e+02| 3.9e+01| 3.1e+02| 4.9e+02
NGC2976_00      |CO10-9 | | 9.8e+01| 1.9e+01| 2.2e+02| 4.0e+02
NGC2976_00      |CO11-10| | 6.4e+01| 7.2e+00| 1.7e+02| 3.9e+02
NGC2976_00      |CO12-11| | 1.2e+02| 3.9e+01| 2.0e+02| 3.6e+02
NGC2976_00      |NII    | | 2.5e+03| 2.4e+03| 2.6e+03|
M81             |CI1-0  | | 1.0e+03| 5.9e+02| 1.4e+03|
M81             |CI2-1  | | 3.1e+02| 2.4e+02| 3.7e+02|
M81             |CO4-3  | | 7.5e+02| 3.4e+02| 1.2e+03| 2.0e+03
M81             |CO5-4  | | 2.4e+02| 4.9e+01| 4.4e+02| 9.8e+02
M81             |CO6-5  | | 2.0e+02| 7.4e+01| 3.2e+02| 4.9e+02
M81             |CO7-6  | | 4.4e+01| 1.2e+01| 1.2e+02| 1.8e+02
M81             |CO8-7  | | 1.1e+02| 4.2e+01| 1.8e+02| 2.4e+02
M81             |CO9-8  | | 1.5e+02| 3.3e+01| 2.8e+02| 4.3e+02
M81             |CO10-9 | | 9.5e+01| 1.6e+01| 1.6e+02| 3.9e+02
M81             |CO12-11| | 1.0e+02| 3.0e+01| 2.2e+02| 4.2e+02
M81             |CO13-12| | 1.8e+02| 4.3e+01| 3.1e+02| 5.3e+02
M81             |NII    | | 2.4e+03| 2.3e+03| 2.6e+03|
M82             |CI1-0  | | 1.7e+04| 1.6e+04| 1.7e+04|
M82             |CI2-1  | | 3.3e+04| 3.2e+04| 3.4e+04|
M82             |CO4-3  | | 5.5e+04| 5.4e+04| 5.6e+04|
M82             |CO5-4  | | 6.3e+04| 6.2e+04| 6.4e+04|
M82             |CO6-5  | | 6.3e+04| 6.2e+04| 6.3e+04|
M82             |CO7-6  | | 5.7e+04| 5.6e+04| 5.8e+04|
M82             |CO8-7  | | 5.1e+04| 5.0e+04| 5.3e+04|
M82             |CO9-8  | | 4.0e+04| 3.9e+04| 4.1e+04|
M82             |CO10-9 | | 3.0e+04| 2.9e+04| 3.0e+04|
M82             |CO11-10| | 2.0e+04| 1.9e+04| 2.0e+04|
M82             |CO12-11| | 1.4e+04| 1.3e+04| 1.5e+04|
M82             |CO13-12| | 8.6e+03| 6.3e+03| 1.1e+04|
M82             |NII    | | 9.0e+04| 8.8e+04| 9.2e+04|
NGC3077         |CI2-1  | | 4.9e+01| 1.4e+01| 9.6e+01| 1.5e+02
NGC3077         |CO4-3  | | 2.2e+02| 7.1e+01| 3.1e+02| 4.8e+02
NGC3077         |CO5-4  | | 1.4e+02| 5.0e+01| 2.6e+02| 4.0e+02
NGC3077         |CO6-5  | | 7.6e+01| 2.4e+01| 1.4e+02| 2.0e+02
NGC3077         |CO7-6  | | 9.2e+01| 4.8e+01| 1.3e+02| 1.9e+02
NGC3077         |CO9-8  | | 3.7e+01| 3.5e+00| 1.0e+02| 2.3e+02
NGC3077         |CO11-10| | 9.8e+01| 2.8e+01| 2.1e+02| 3.5e+02
NGC3077         |CO12-11| | 7.7e+01| 1.8e+01| 1.6e+02| 2.7e+02
NGC3077         |CO13-12| | 1.5e+02| 6.0e+01| 2.6e+02| 4.6e+02
NGC3077         |NII    | | 3.8e+03| 3.6e+03| 3.9e+03|
NGC3110a        |CI1-0  | | 9.9e+02| 4.8e+02| 1.4e+03| 2.1e+03
NGC3110a        |CI2-1  | | 7.3e+02| 6.1e+02| 8.3e+02|
NGC3110a        |CO5-4  | | 4.9e+02| 1.8e+02| 8.6e+02| 1.6e+03
NGC3110a        |CO6-5  | | 5.9e+02| 3.2e+02| 7.8e+02|
NGC3110a        |CO7-6  | | 4.0e+02| 2.7e+02| 5.0e+02|
NGC3110a        |CO8-7  | | 1.8e+02| 5.6e+01| 3.4e+02| 5.7e+02
NGC3110a        |CO9-8  | | 3.7e+02| 1.7e+02| 5.7e+02| 8.3e+02
NGC3110a        |CO10-9 | | 2.3e+02| 8.1e+01| 3.7e+02| 5.4e+02
NGC3110a        |CO12-11| | 1.4e+02| 3.9e+01| 2.7e+02| 4.6e+02
NGC3110a        |NII    | | 3.1e+03| 3.0e+03| 3.2e+03|
3C 236          |CO5-4  | | 1.7e+02| 4.7e+01| 2.9e+02| 4.9e+02
3C 236          |CO6-5  | | 6.6e+01| 2.4e+01| 1.1e+02| 1.8e+02
3C 236          |CO8-7  | | 5.9e+01| 2.0e+01| 9.9e+01| 1.6e+02
3C 236          |CO11-10| | 2.0e+01| 2.9e+00| 4.7e+01| 8.9e+01
3C 236          |CO12-11| | 3.5e+01| 1.0e+01| 7.2e+01| 1.2e+02
3C 236          |NII    | | 2.8e+01| 1.0e+01| 6.7e+01| 1.2e+02
NGC3221         |CI1-0  | | 3.5e+02| 1.0e+02| 7.9e+02| 1.0e+03
NGC3221         |CI2-1  | | 3.7e+02| 2.2e+02| 4.9e+02|
NGC3221         |CO4-3  | | 7.1e+02| 2.6e+02| 1.1e+03| 1.6e+03
NGC3221         |CO5-4  | | 5.8e+02| 2.7e+02| 9.1e+02| 1.4e+03
NGC3221         |CO6-5  | | 2.8e+02| 1.1e+02| 4.6e+02| 7.5e+02
NGC3221         |CO8-7  | | 1.2e+02| 2.0e+01| 2.8e+02| 5.6e+02
NGC3221         |CO9-8  | | 4.4e+02| 1.2e+02| 7.3e+02| 1.2e+03
NGC3221         |CO10-9 | | 3.8e+02| 1.2e+02| 6.9e+02| 1.0e+03
NGC3221         |CO12-11| | 2.4e+02| 5.6e+01| 4.2e+02| 6.9e+02
NGC3221         |NII    | | 3.4e+03| 3.1e+03| 3.7e+03|
NGC3227         |CI1-0  | | 1.1e+03| 8.6e+02| 1.4e+03|
NGC3227         |CI2-1  | | 1.8e+03| 1.7e+03| 1.8e+03|
NGC3227         |CO4-3  | | 1.7e+03| 1.4e+03| 2.0e+03|
NGC3227         |CO5-4  | | 1.6e+03| 1.4e+03| 1.8e+03|
NGC3227         |CO6-5  | | 1.2e+03| 1.1e+03| 1.3e+03|
NGC3227         |CO7-6  | | 7.4e+02| 6.7e+02| 8.0e+02|
NGC3227         |CO8-7  | | 7.0e+02| 6.1e+02| 7.9e+02|
NGC3227         |CO9-8  | | 4.4e+02| 3.1e+02| 5.8e+02|
NGC3227         |CO10-9 | | 3.3e+02| 2.0e+02| 4.3e+02|
NGC3227         |CO11-10| | 4.0e+02| 2.7e+02| 5.1e+02|
NGC3227         |CO12-11| | 3.1e+02| 2.2e+02| 4.0e+02|
NGC3227         |CO13-12| | 1.0e+02| 2.8e+01| 1.9e+02| 3.5e+02
NGC3227         |NII    |X| 2.0e+03| 1.9e+03| 2.2e+03|
NGC3256         |CI1-0  | | 3.3e+03| 3.1e+03| 3.6e+03|
NGC3256         |CI2-1  | | 4.8e+03| 4.7e+03| 4.9e+03|
NGC3256         |CO4-3  | | 8.4e+03| 8.2e+03| 8.8e+03|
NGC3256         |CO5-4  | | 8.3e+03| 8.1e+03| 8.4e+03|
NGC3256         |CO6-5  | | 8.2e+03| 8.2e+03| 8.4e+03|
NGC3256         |CO7-6  | | 5.7e+03| 5.6e+03| 5.8e+03|
NGC3256         |CO8-7  | | 4.4e+03| 4.2e+03| 4.5e+03|
NGC3256         |CO9-8  | | 3.1e+03| 2.9e+03| 3.2e+03|
NGC3256         |CO10-9 | | 2.2e+03| 2.0e+03| 2.3e+03|
NGC3256         |CO11-10| | 1.4e+03| 1.2e+03| 1.4e+03|
NGC3256         |CO12-11| | 9.2e+02| 8.2e+02| 1.0e+03|
NGC3256         |CO13-12| | 5.2e+02| 2.9e+02| 7.2e+02|
NGC3256         |NII    | | 9.3e+03| 9.1e+03| 9.5e+03|
IRAS 10378+1109 |CI2-1  | | 6.2e+01| 2.4e+01| 1.0e+02| 1.6e+02
IRAS 10378+1109 |CO5-4  | | 1.0e+02| 3.8e+01| 2.1e+02| 3.8e+02
IRAS 10378+1109 |CO6-5  | | 1.7e+02| 7.3e+01| 2.4e+02| 3.5e+02
IRAS 10378+1109 |CO7-6  | | 2.2e+02| 1.8e+02| 2.5e+02|
IRAS 10378+1109 |CO8-7  | | 1.5e+02| 1.1e+02| 1.8e+02|
IRAS 10378+1109 |CO10-9 | | 9.2e+01| 5.5e+01| 1.4e+02| 2.0e+02
IRAS 10378+1109 |CO11-10| | 3.2e+01| 8.5e+00| 5.6e+01| 1.1e+02
IRAS 10378+1109 |CO12-11| | 2.1e+01| 3.7e+00| 4.4e+01| 8.2e+01
IRAS 10378+1109 |CO13-12| | 7.1e+01| 4.8e+01| 1.0e+02| 1.5e+02
IRAS 10378+1109 |NII    | | 7.0e+01| 4.4e+01| 1.0e+02| 1.5e+02
ESO264-G036     |CI1-0  | | 4.6e+02| 1.9e+02| 6.8e+02| 9.7e+02
ESO264-G036     |CI2-1  | | 4.9e+02| 4.4e+02| 5.4e+02|
ESO264-G036     |CO5-4  | | 6.2e+02| 4.7e+02| 7.4e+02|
ESO264-G036     |CO6-5  | | 5.8e+02| 4.9e+02| 6.6e+02|
ESO264-G036     |CO7-6  | | 3.1e+02| 2.6e+02| 3.6e+02|
ESO264-G036     |CO8-7  | | 3.1e+02| 2.2e+02| 3.9e+02|
ESO264-G036     |CO9-8  | | 1.0e+02| 2.9e+01| 2.0e+02| 3.6e+02
ESO264-G036     |CO10-9 | | 1.2e+02| 4.1e+01| 2.2e+02| 3.6e+02
ESO264-G036     |CO12-11| | 9.2e+01| 2.9e+01| 2.0e+02| 3.1e+02
ESO264-G036     |NII    |X| 3.2e+03| 3.1e+03| 3.3e+03|
NGC3351         |CI1-0  | | 6.7e+02| 4.6e+02| 9.0e+02|
NGC3351         |CI2-1  | | 6.8e+02| 6.2e+02| 7.4e+02|
NGC3351         |CO4-3  | | 1.0e+03| 8.4e+02| 1.3e+03|
NGC3351         |CO5-4  | | 1.2e+03| 1.1e+03| 1.4e+03|
NGC3351         |CO6-5  | | 6.7e+02| 5.8e+02| 7.6e+02|
NGC3351         |CO7-6  | | 3.8e+02| 3.2e+02| 4.4e+02|
NGC3351         |CO8-7  | | 1.8e+02| 1.1e+02| 2.6e+02| 3.4e+02
NGC3351         |CO9-8  | | 3.2e+02| 2.0e+02| 4.6e+02|
NGC3351         |CO10-9 | | 1.8e+02| 9.1e+01| 2.8e+02| 4.2e+02
NGC3351         |CO11-10| | 1.2e+02| 3.4e+01| 2.2e+02| 4.3e+02
NGC3351         |CO12-11| | 1.2e+02| 3.2e+01| 2.1e+02| 3.3e+02
NGC3351         |CO13-12| | 3.6e+02| 2.2e+02| 5.2e+02|
NGC3351         |NII    | | 6.5e+03| 6.4e+03| 6.6e+03|
ESO264-G057     |CI1-0  | | 2.5e+02| 1.0e+02| 4.2e+02| 6.6e+02
ESO264-G057     |CI2-1  | | 2.4e+02| 2.0e+02| 3.0e+02|
ESO264-G057     |CO5-4  | | 2.8e+02| 1.6e+02| 3.9e+02|
ESO264-G057     |CO6-5  | | 3.0e+02| 2.4e+02| 3.7e+02|
ESO264-G057     |CO7-6  | | 2.0e+02| 1.5e+02| 2.5e+02|
ESO264-G057     |CO8-7  | | 2.4e+02| 1.5e+02| 3.2e+02|
ESO264-G057     |CO9-8  | | 1.0e+02| 2.3e+01| 1.8e+02| 3.7e+02
ESO264-G057     |CO10-9 | | 1.5e+02| 4.9e+01| 2.3e+02| 3.4e+02
ESO264-G057     |CO11-10| | 1.2e+02| 4.2e+01| 2.0e+02| 3.6e+02
ESO264-G057     |CO12-11| | 6.9e+01| 1.8e+01| 1.8e+02| 2.8e+02
ESO264-G057     |NII    | | 1.7e+03| 1.6e+03| 1.8e+03|
IRASF10565+2448 |CI1-0  | | 3.6e+02| 8.7e+01| 7.1e+02| 1.1e+03
IRASF10565+2448 |CI2-1  | | 5.2e+02| 4.5e+02| 5.8e+02|
IRASF10565+2448 |CO5-4  | | 6.4e+02| 4.3e+02| 8.2e+02|
IRASF10565+2448 |CO6-5  | | 7.5e+02| 6.6e+02| 8.3e+02|
IRASF10565+2448 |CO7-6  | | 5.4e+02| 4.7e+02| 6.1e+02|
IRASF10565+2448 |CO8-7  | | 6.1e+02| 5.4e+02| 6.9e+02|
IRASF10565+2448 |CO9-8  | | 3.8e+02| 3.0e+02| 4.7e+02|
IRASF10565+2448 |CO10-9 | | 3.2e+02| 2.6e+02| 3.9e+02|
IRASF10565+2448 |CO11-10| | 2.4e+02| 1.8e+02| 3.0e+02|
IRASF10565+2448 |CO12-11| | 1.2e+02| 6.5e+01| 1.7e+02|
IRASF10565+2448 |CO13-12| | 9.3e+01| 3.9e+01| 1.4e+02| 2.2e+02
IRASF10565+2448 |NII    | | 5.0e+02| 4.6e+02| 5.5e+02|
NGC3521         |CI1-0  | | 1.3e+03| 1.0e+03| 1.5e+03|
NGC3521         |CI2-1  | | 9.2e+02| 8.3e+02| 1.0e+03|
NGC3521         |CO4-3  | | 1.5e+03| 1.3e+03| 1.8e+03|
NGC3521         |CO5-4  | | 7.5e+02| 5.5e+02| 1.0e+03|
NGC3521         |CO6-5  | | 3.0e+02| 1.8e+02| 4.2e+02|
NGC3521         |CO7-6  | | 6.1e+01| 1.2e+01| 1.2e+02| 2.2e+02
NGC3521         |CO9-8  | | 1.9e+02| 3.6e+01| 4.3e+02| 1.0e+03
NGC3521         |CO12-11| | 4.8e+02| 1.8e+02| 7.3e+02| 1.1e+03
NGC3521         |NII    | | 1.1e+04| 1.1e+04| 1.1e+04|
IRAS 11095-0238 |CO5-4  | | 1.5e+02| 4.1e+01| 2.7e+02| 4.1e+02
IRAS 11095-0238 |CO6-5  | | 6.9e+01| 1.8e+01| 1.1e+02| 1.6e+02
IRAS 11095-0238 |CO7-6  | | 1.3e+02| 7.6e+01| 1.7e+02|
IRAS 11095-0238 |CO8-7  | | 1.6e+02| 1.1e+02| 2.0e+02|
IRAS 11095-0238 |CO10-9 | | 1.3e+02| 8.0e+01| 1.8e+02|
IRAS 11095-0238 |CO11-10| | 6.0e+01| 2.4e+01| 1.1e+02| 1.6e+02
IRAS 11095-0238 |CO12-11| | 6.7e+01| 2.2e+01| 1.1e+02| 1.6e+02
IRAS 11095-0238 |CO13-12| | 5.8e+01| 2.8e+01| 9.3e+01| 1.5e+02
IRAS 11095-0238 |NII    | | 1.0e+02| 6.7e+01| 1.3e+02|
NGC3627         |CI1-0  | | 1.4e+03| 1.3e+03| 1.6e+03|
NGC3627         |CI2-1  | | 1.2e+03| 1.1e+03| 1.2e+03|
NGC3627         |CO4-3  | | 1.6e+03| 1.4e+03| 1.8e+03|
NGC3627         |CO5-4  | | 2.4e+03| 2.2e+03| 2.5e+03|
NGC3627         |CO6-5  | | 2.0e+03| 1.9e+03| 2.0e+03|
NGC3627         |CO7-6  | | 1.3e+03| 1.2e+03| 1.3e+03|
NGC3627         |CO8-7  | | 9.3e+02| 8.6e+02| 9.9e+02|
NGC3627         |CO9-8  | | 1.4e+03| 1.2e+03| 1.5e+03|
NGC3627         |CO10-9 | | 1.2e+03| 1.1e+03| 1.3e+03|
NGC3627         |CO11-10| | 6.3e+02| 5.0e+02| 7.6e+02|
NGC3627         |CO12-11| | 3.7e+02| 2.7e+02| 4.7e+02|
NGC3627         |CO13-12| | 3.6e+02| 1.7e+02| 5.4e+02|
NGC3627         |NII    | | 1.9e+03| 1.7e+03| 2.0e+03|
NGC3665         |CI1-0  | | 1.3e+02| 3.8e+01| 2.4e+02| 4.5e+02
NGC3665         |CI2-1  | | 1.2e+02| 9.4e+01| 1.5e+02|
NGC3665         |CO4-3  | | 2.1e+02| 6.2e+01| 3.8e+02| 5.6e+02
NGC3665         |CO5-4  | | 8.5e+01| 2.5e+01| 1.7e+02| 2.7e+02
NGC3665         |CO6-5  | | 6.4e+01| 2.5e+01| 1.0e+02| 1.5e+02
NGC3665         |CO7-6  | | 1.7e+01| 2.9e+00| 3.8e+01| 6.1e+01
NGC3665         |CO8-7  | | 6.8e+01| 2.4e+01| 1.2e+02| 1.8e+02
NGC3665         |CO9-8  | | 5.6e+01| 1.7e+01| 9.2e+01| 1.6e+02
NGC3665         |NII    |X| 1.5e+03| 1.4e+03| 1.5e+03|
Arp299-B        |CI1-0  | | 2.1e+03| 1.6e+03| 2.5e+03|
Arp299-B        |CI2-1  | | 2.1e+03| 2.0e+03| 2.2e+03|
Arp299-B        |CO4-3  | | 5.9e+03| 5.4e+03| 6.3e+03|
Arp299-B        |CO5-4  | | 5.2e+03| 4.9e+03| 5.5e+03|
Arp299-B        |CO6-5  | | 4.5e+03| 4.4e+03| 4.7e+03|
Arp299-B        |CO7-6  | | 3.1e+03| 3.0e+03| 3.2e+03|
Arp299-B        |CO8-7  | | 2.6e+03| 2.5e+03| 2.8e+03|
Arp299-B        |CO9-8  | | 1.7e+03| 1.4e+03| 1.9e+03|
Arp299-B        |CO10-9 | | 1.6e+03| 1.4e+03| 1.8e+03|
Arp299-B        |CO11-10| | 1.4e+03| 1.2e+03| 1.5e+03|
Arp299-B        |CO12-11| | 1.1e+03| 9.7e+02| 1.3e+03|
Arp299-B        |CO13-12| | 1.0e+03| 8.3e+02| 1.2e+03|
Arp299-B        |NII    |X| 8.2e+03| 7.9e+03| 8.5e+03|
Arp299-C        |CI1-0  | | 2.0e+03| 1.6e+03| 2.4e+03|
Arp299-C        |CI2-1  | | 2.0e+03| 1.9e+03| 2.1e+03|
Arp299-C        |CO4-3  | | 5.7e+03| 5.2e+03| 6.1e+03|
Arp299-C        |CO5-4  | | 5.6e+03| 5.4e+03| 5.9e+03|
Arp299-C        |CO6-5  | | 4.2e+03| 4.0e+03| 4.4e+03|
Arp299-C        |CO7-6  | | 3.0e+03| 2.9e+03| 3.1e+03|
Arp299-C        |CO8-7  | | 2.7e+03| 2.6e+03| 2.9e+03|
Arp299-C        |CO9-8  | | 1.7e+03| 1.5e+03| 1.8e+03|
Arp299-C        |CO10-9 | | 1.4e+03| 1.2e+03| 1.5e+03|
Arp299-C        |CO11-10| | 1.1e+03| 9.8e+02| 1.3e+03|
Arp299-C        |CO12-11| | 7.7e+02| 6.3e+02| 9.1e+02|
Arp299-C        |CO13-12| | 5.0e+02| 3.3e+02| 6.8e+02|
Arp299-C        |NII    |X| 7.7e+03| 7.4e+03| 7.9e+03|
Arp299-A        |CI1-0  | | 1.3e+03| 1.1e+03| 1.6e+03|
Arp299-A        |CI2-1  | | 2.3e+03| 2.2e+03| 2.4e+03|
Arp299-A        |CO4-3  | | 5.1e+03| 4.8e+03| 5.4e+03|
Arp299-A        |CO5-4  | | 4.8e+03| 4.7e+03| 5.0e+03|
Arp299-A        |CO6-5  | | 4.7e+03| 4.6e+03| 4.8e+03|
Arp299-A        |CO7-6  | | 4.0e+03| 3.9e+03| 4.1e+03|
Arp299-A        |CO8-7  | | 3.7e+03| 3.6e+03| 3.8e+03|
Arp299-A        |CO9-8  | | 3.2e+03| 3.0e+03| 3.3e+03|
Arp299-A        |CO10-9 | | 2.9e+03| 2.7e+03| 3.0e+03|
Arp299-A        |CO11-10| | 2.2e+03| 2.1e+03| 2.4e+03|
Arp299-A        |CO12-11| | 1.8e+03| 1.7e+03| 1.9e+03|
Arp299-A        |CO13-12| | 1.6e+03| 1.4e+03| 1.7e+03|
Arp299-A        |NII    |X| 5.6e+03| 5.3e+03| 5.8e+03|
PG 1126-041     |CI2-1  | | 3.0e+01| 4.4e+00| 6.7e+01| 9.7e+01
PG 1126-041     |CO6-5  | | 6.6e+01| 2.2e+01| 1.1e+02| 2.0e+02
PG 1126-041     |CO7-6  | | 2.8e+01| 4.8e+00| 6.1e+01| 1.1e+02
PG 1126-041     |CO8-7  | | 2.3e+01| 4.5e+00| 5.8e+01| 9.8e+01
PG 1126-041     |CO9-8  | | 9.4e+01| 5.2e+01| 1.4e+02| 2.4e+02
PG 1126-041     |CO10-9 | | 4.4e+01| 1.6e+01| 7.6e+01| 1.3e+02
PG 1126-041     |CO11-10| | 5.4e+01| 2.3e+01| 8.4e+01| 1.3e+02
PG 1126-041     |CO12-11| | 6.9e+01| 3.5e+01| 1.0e+02| 1.5e+02
PG 1126-041     |CO13-12| | 2.4e+01| 4.8e+00| 6.0e+01| 9.0e+01
PG 1126-041     |NII    | | 9.4e+01| 6.7e+01| 1.3e+02|
ESO 320-G030    |CI1-0  | | 9.4e+02| 6.9e+02| 1.2e+03|
ESO 320-G030    |CI2-1  | | 8.5e+02| 7.8e+02| 9.1e+02|
ESO 320-G030    |CO4-3  | | 2.6e+03| 2.3e+03| 2.8e+03|
ESO 320-G030    |CO5-4  | | 2.0e+03| 1.8e+03| 2.1e+03|
ESO 320-G030    |CO6-5  | | 1.8e+03| 1.7e+03| 1.9e+03|
ESO 320-G030    |CO7-6  | | 1.2e+03| 1.2e+03| 1.3e+03|
ESO 320-G030    |CO8-7  | | 8.1e+02| 7.3e+02| 8.9e+02|
ESO 320-G030    |CO9-8  | | 8.0e+02| 7.0e+02| 8.9e+02|
ESO 320-G030    |CO10-9 | | 7.6e+02| 6.8e+02| 8.3e+02|
ESO 320-G030    |CO11-10| | 3.4e+02| 2.7e+02| 4.2e+02|
ESO 320-G030    |CO12-11| | 2.6e+02| 2.0e+02| 3.1e+02|
ESO 320-G030    |CO13-12| | 1.4e+02| 5.7e+01| 2.0e+02| 3.5e+02
ESO 320-G030    |NII    | | 2.3e+03| 2.2e+03| 2.4e+03|
NGC3982         |CI1-0  | | 5.8e+02| 2.7e+02| 7.9e+02|
NGC3982         |CI2-1  | | 3.9e+02| 3.4e+02| 4.5e+02|
NGC3982         |CO4-3  | | 1.1e+03| 7.2e+02| 1.4e+03|
NGC3982         |CO5-4  | | 3.4e+02| 1.7e+02| 5.1e+02| 8.2e+02
NGC3982         |CO6-5  | | 3.4e+02| 2.4e+02| 4.5e+02|
NGC3982         |CO7-6  | | 1.2e+02| 4.6e+01| 1.8e+02| 2.8e+02
NGC3982         |CO8-7  | | 9.9e+01| 2.5e+01| 1.7e+02| 3.2e+02
NGC3982         |CO9-8  | | 6.0e+01| 5.7e+00| 1.5e+02| 3.5e+02
NGC3982         |CO11-10| | 2.6e+02| 8.7e+01| 4.3e+02| 6.0e+02
NGC3982         |NII    | | 4.4e+03| 4.3e+03| 4.6e+03|
NGC4038         |CI1-0  | | 3.8e+02| 1.8e+02| 6.4e+02| 8.4e+02
NGC4038         |CI2-1  | | 9.8e+02| 8.6e+02| 1.1e+03|
NGC4038         |CO4-3  | | 1.2e+03| 8.8e+02| 1.4e+03|
NGC4038         |CO5-4  | | 1.2e+03| 9.0e+02| 1.5e+03|
NGC4038         |CO6-5  | | 1.2e+03| 1.0e+03| 1.3e+03|
NGC4038         |CO7-6  | | 9.0e+02| 7.5e+02| 1.0e+03|
NGC4038         |CO8-7  | | 2.8e+02| 9.3e+01| 4.6e+02| 7.3e+02
NGC4038         |CO9-8  | | 5.2e+02| 2.5e+02| 8.8e+02| 1.4e+03
NGC4038         |CO12-11| | 1.7e+02| 2.2e+01| 3.5e+02| 5.9e+02
NGC4038         |CO13-12| | 5.4e+02| 2.0e+02| 8.3e+02| 1.2e+03
NGC4038         |NII    | | 3.2e+03| 2.9e+03| 3.4e+03|
NGC4038overlap  |CI1-0  | | 6.7e+02| 3.4e+02| 1.0e+03|
NGC4038overlap  |CI2-1  | | 1.5e+03| 1.4e+03| 1.6e+03|
NGC4038overlap  |CO4-3  | | 2.4e+03| 1.9e+03| 2.8e+03|
NGC4038overlap  |CO5-4  | | 2.0e+03| 1.8e+03| 2.3e+03|
NGC4038overlap  |CO6-5  | | 1.8e+03| 1.6e+03| 1.9e+03|
NGC4038overlap  |CO7-6  | | 1.3e+03| 1.2e+03| 1.4e+03|
NGC4038overlap  |CO8-7  | | 9.4e+02| 7.6e+02| 1.1e+03|
NGC4038overlap  |CO9-8  | | 2.6e+02| 7.8e+01| 5.3e+02| 1.0e+03
NGC4038overlap  |CO10-9 | | 5.8e+02| 2.7e+02| 8.6e+02| 1.3e+03
NGC4038overlap  |CO12-11| | 4.5e+02| 1.7e+02| 7.1e+02| 1.1e+03
NGC4038overlap  |CO13-12| | 4.2e+02| 1.4e+02| 7.8e+02| 1.3e+03
NGC4038overlap  |NII    | | 4.2e+03| 3.9e+03| 4.5e+03|
NGC4051         |CI1-0  | | 7.4e+02| 4.8e+02| 1.0e+03|
NGC4051         |CI2-1  | | 5.3e+02| 4.6e+02| 6.0e+02|
NGC4051         |CO4-3  | | 8.2e+02| 5.0e+02| 1.1e+03| 1.6e+03
NGC4051         |CO5-4  | | 6.1e+02| 4.1e+02| 8.1e+02|
NGC4051         |CO6-5  | | 6.8e+02| 5.9e+02| 7.7e+02|
NGC4051         |CO7-6  | | 4.1e+02| 3.3e+02| 4.9e+02|
NGC4051         |CO8-7  | | 4.4e+02| 3.5e+02| 5.4e+02|
NGC4051         |CO9-8  | | 4.4e+02| 2.8e+02| 6.0e+02|
NGC4051         |CO10-9 | | 1.4e+02| 3.9e+01| 2.6e+02| 4.9e+02
NGC4051         |CO11-10| | 3.0e+02| 1.9e+02| 4.4e+02|
NGC4051         |CO12-11| | 1.1e+02| 3.0e+01| 1.9e+02| 3.6e+02
NGC4051         |CO13-12| | 2.3e+02| 9.8e+01| 3.5e+02| 5.2e+02
NGC4051         |NII    | | 8.4e+02| 7.2e+02| 9.3e+02|
IRAS 12071-0444 |CI2-1  | | 6.3e+01| 2.5e+01| 9.9e+01| 1.5e+02
IRAS 12071-0444 |CO5-4  | | 2.1e+02| 1.0e+02| 3.3e+02| 5.6e+02
IRAS 12071-0444 |CO6-5  | | 1.5e+02| 8.6e+01| 2.2e+02| 3.6e+02
IRAS 12071-0444 |CO7-6  | | 9.0e+01| 4.8e+01| 1.3e+02|
IRAS 12071-0444 |CO8-7  | | 1.4e+02| 1.0e+02| 1.7e+02|
IRAS 12071-0444 |CO10-9 | | 9.2e+01| 4.3e+01| 1.4e+02| 2.2e+02
IRAS 12071-0444 |CO11-10| | 4.6e+01| 1.6e+01| 8.2e+01| 1.4e+02
IRAS 12071-0444 |CO12-11| | 7.3e+01| 3.7e+01| 1.1e+02| 1.5e+02
IRAS 12071-0444 |CO13-12| | 4.0e+01| 1.4e+01| 6.8e+01| 1.2e+02
IRAS 12071-0444 |NII    | | 4.9e+01| 2.0e+01| 8.1e+01| 1.4e+02
NGC4151         |CI1-0  | | 2.8e+02| 1.1e+02| 5.3e+02| 8.5e+02
NGC4151         |CI2-1  | | 4.8e+02| 4.3e+02| 5.5e+02|
NGC4151         |CO4-3  | | 2.2e+02| 6.8e+01| 4.6e+02| 8.9e+02
NGC4151         |CO6-5  | | 1.1e+02| 4.4e+01| 1.8e+02| 3.0e+02
NGC4151         |CO7-6  | | 1.7e+02| 1.1e+02| 2.3e+02|
NGC4151         |CO8-7  | | 1.8e+02| 1.1e+02| 2.4e+02| 3.4e+02
NGC4151         |CO9-8  | | 1.9e+02| 8.6e+01| 2.8e+02| 4.0e+02
NGC4151         |CO10-9 | | 4.7e+02| 3.7e+02| 5.8e+02|
NGC4151         |CO11-10| | 1.6e+02| 8.8e+01| 2.6e+02| 4.1e+02
NGC4151         |CO12-11| | 1.1e+02| 3.3e+01| 1.8e+02| 3.2e+02
NGC4151         |CO13-12| | 2.1e+02| 1.2e+02| 3.1e+02|
NGC4151         |NII    |X| 1.4e+03| 1.2e+03| 1.5e+03|
NGC4194         |CI1-0  | | 5.0e+02| 2.3e+02| 8.7e+02| 1.4e+03
NGC4194         |CI2-1  | | 5.4e+02| 4.4e+02| 6.1e+02|
NGC4194         |CO4-3  | | 8.3e+02| 4.9e+02| 1.2e+03|
NGC4194         |CO5-4  | | 5.0e+02| 2.2e+02| 7.0e+02|
NGC4194         |CO6-5  | | 9.1e+02| 8.0e+02| 1.0e+03|
NGC4194         |CO7-6  | | 9.0e+02| 8.2e+02| 9.7e+02|
NGC4194         |CO8-7  | | 5.6e+02| 4.4e+02| 6.9e+02|
NGC4194         |CO9-8  | | 2.8e+02| 1.1e+02| 4.4e+02| 6.7e+02
NGC4194         |CO10-9 | | 3.0e+02| 1.6e+02| 4.2e+02|
NGC4194         |CO11-10| | 5.2e+02| 4.0e+02| 6.5e+02|
NGC4194         |CO12-11| | 2.7e+02| 1.8e+02| 3.6e+02|
NGC4194         |CO13-12| | 1.9e+02| 7.5e+01| 2.9e+02| 4.5e+02
NGC4194         |NII    | | 1.7e+03| 1.6e+03| 1.8e+03|
IRAS12116-5615  |CI1-0  | | 3.9e+02| 1.8e+02| 5.9e+02| 9.8e+02
IRAS12116-5615  |CI2-1  | | 5.6e+02| 5.1e+02| 6.2e+02|
IRAS12116-5615  |CO5-4  | | 8.1e+02| 6.4e+02| 9.4e+02|
IRAS12116-5615  |CO6-5  | | 6.9e+02| 6.1e+02| 7.6e+02|
IRAS12116-5615  |CO7-6  | | 5.8e+02| 5.2e+02| 6.3e+02|
IRAS12116-5615  |CO8-7  | | 4.3e+02| 3.6e+02| 4.9e+02|
IRAS12116-5615  |CO9-8  | | 4.0e+02| 3.2e+02| 4.8e+02|
IRAS12116-5615  |CO10-9 | | 2.0e+02| 1.4e+02| 2.6e+02|
IRAS12116-5615  |CO11-10| | 1.5e+02| 9.0e+01| 2.0e+02|
IRAS12116-5615  |CO12-11| | 1.0e+02| 4.7e+01| 1.5e+02|
IRAS12116-5615  |CO13-12| | 9.3e+01| 4.0e+01| 1.4e+02| 2.1e+02
IRAS12116-5615  |NII    | | 7.1e+02| 6.6e+02| 7.5e+02|
NGC4254         |CI1-0  | | 1.0e+03| 8.6e+02| 1.2e+03|
NGC4254         |CI2-1  | | 6.8e+02| 6.2e+02| 7.5e+02|
NGC4254         |CO4-3  | | 6.4e+02| 4.3e+02| 8.9e+02|
NGC4254         |CO5-4  | | 5.9e+02| 3.6e+02| 8.0e+02|
NGC4254         |CO6-5  | | 2.0e+02| 8.7e+01| 2.9e+02| 4.3e+02
NGC4254         |CO7-6  | | 7.2e+01| 1.4e+01| 1.4e+02| 2.4e+02
NGC4254         |CO9-8  | | 2.2e+02| 4.8e+01| 3.9e+02| 6.0e+02
NGC4254         |CO11-10| | 1.5e+02| 2.3e+01| 3.3e+02| 6.2e+02
NGC4254         |NII    | | 1.2e+04| 1.2e+04| 1.2e+04|
NGC4321         |CI1-0  | | 1.0e+03| 8.6e+02| 1.2e+03|
NGC4321         |CI2-1  | | 8.5e+02| 8.0e+02| 9.0e+02|
NGC4321         |CO4-3  | | 2.4e+03| 2.2e+03| 2.6e+03|
NGC4321         |CO5-4  | | 1.7e+03| 1.6e+03| 1.9e+03|
NGC4321         |CO6-5  | | 1.2e+03| 1.1e+03| 1.3e+03|
NGC4321         |CO7-6  | | 5.3e+02| 4.8e+02| 5.8e+02|
NGC4321         |CO8-7  | | 1.9e+02| 1.0e+02| 2.8e+02| 3.5e+02
NGC4321         |CO9-8  | | 1.0e+02| 2.5e+01| 2.4e+02| 3.9e+02
NGC4321         |CO10-9 | | 3.7e+02| 2.4e+02| 4.6e+02|
NGC4321         |CO11-10| | 3.2e+02| 1.8e+02| 4.5e+02| 6.2e+02
NGC4321         |CO13-12| | 2.4e+02| 7.7e+01| 4.2e+02| 6.8e+02
NGC4321         |NII    | | 8.9e+03| 8.7e+03| 9.0e+03|
NGC4388         |CI1-0  | | 9.2e+02| 6.3e+02| 1.2e+03|
NGC4388         |CI2-1  | | 1.2e+03| 1.1e+03| 1.2e+03|
NGC4388         |CO4-3  | | 1.6e+03| 1.3e+03| 1.9e+03|
NGC4388         |CO5-4  | | 9.5e+02| 7.6e+02| 1.1e+03|
NGC4388         |CO6-5  | | 8.5e+02| 7.5e+02| 9.4e+02|
NGC4388         |CO7-6  | | 5.7e+02| 5.2e+02| 6.2e+02|
NGC4388         |CO8-7  | | 4.9e+02| 4.0e+02| 5.6e+02|
NGC4388         |CO9-8  | | 3.9e+02| 2.4e+02| 5.3e+02|
NGC4388         |CO10-9 | | 2.9e+02| 2.0e+02| 4.2e+02|
NGC4388         |CO11-10| | 1.7e+02| 7.3e+01| 3.1e+02| 4.8e+02
NGC4388         |CO12-11| | 1.5e+02| 5.7e+01| 2.5e+02| 4.1e+02
NGC4388         |CO13-12| | 1.1e+02| 3.7e+01| 2.1e+02| 3.6e+02
NGC4388         |NII    | | 1.9e+03| 1.8e+03| 2.0e+03|
NGC4459         |CI1-0  | | 3.0e+02| 9.2e+01| 6.2e+02| 9.9e+02
NGC4459         |CI2-1  | | 2.3e+02| 1.4e+02| 3.0e+02|
NGC4459         |CO4-3  | | 4.1e+02| 1.3e+02| 7.8e+02| 1.2e+03
NGC4459         |CO5-4  | | 1.4e+02| 2.1e+01| 3.2e+02| 5.9e+02
NGC4459         |CO6-5  | | 3.0e+02| 2.0e+02| 4.2e+02|
NGC4459         |CO9-8  | | 4.4e+01| 1.2e+01| 9.1e+01| 1.6e+02
NGC4459         |CO10-9 | | 6.1e+01| 2.2e+01| 1.0e+02| 1.7e+02
NGC4459         |CO12-11| | 3.8e+01| 1.1e+01| 6.7e+01| 1.2e+02
NGC4459         |CO13-12| | 2.8e+01| 7.1e+00| 6.2e+01| 1.0e+02
NGC4459         |NII    |X| 7.8e+02| 7.4e+02| 8.4e+02|
NGC4526         |CI1-0  | | 4.8e+02| 2.7e+02| 6.2e+02|
NGC4526         |CI2-1  | | 2.2e+02| 1.8e+02| 2.5e+02|
NGC4526         |CO4-3  | | 6.7e+02| 4.5e+02| 8.6e+02|
NGC4526         |CO5-4  | | 3.4e+02| 2.3e+02| 4.3e+02|
NGC4526         |CO6-5  | | 1.9e+02| 1.4e+02| 2.4e+02|
NGC4526         |CO7-6  | | 4.7e+01| 1.9e+01| 8.0e+01| 1.3e+02
NGC4526         |CO8-7  | | 5.4e+01| 1.2e+01| 9.6e+01| 1.8e+02
NGC4526         |CO9-8  | | 4.5e+01| 1.4e+01| 8.4e+01| 1.7e+02
NGC4526         |CO10-9 | | 4.6e+01| 1.5e+01| 8.5e+01| 1.6e+02
NGC4526         |CO12-11| | 5.8e+01| 2.5e+01| 9.4e+01| 1.4e+02
NGC4526         |CO13-12| | 6.4e+01| 2.1e+01| 1.2e+02| 2.1e+02
NGC4526         |NII    |X| 5.3e+03| 5.2e+03| 5.4e+03|
NGC4536         |CI1-0  | | 2.0e+02| 4.6e+01| 4.7e+02| 8.6e+02
NGC4536         |CI2-1  | | 8.8e+02| 8.0e+02| 9.6e+02|
NGC4536         |CO4-3  | | 1.6e+03| 1.3e+03| 2.0e+03|
NGC4536         |CO5-4  | | 1.3e+03| 1.0e+03| 1.5e+03|
NGC4536         |CO6-5  | | 1.3e+03| 1.2e+03| 1.4e+03|
NGC4536         |CO7-6  | | 7.9e+02| 7.0e+02| 8.7e+02|
NGC4536         |CO8-7  | | 4.4e+02| 3.4e+02| 5.5e+02|
NGC4536         |CO9-8  | | 4.5e+02| 2.9e+02| 6.1e+02| 8.3e+02
NGC4536         |CO10-9 | | 3.7e+02| 1.9e+02| 5.0e+02|
NGC4536         |CO11-10| | 2.4e+02| 9.2e+01| 3.9e+02| 5.7e+02
NGC4536         |CO12-11| | 1.3e+02| 2.8e+01| 2.6e+02| 4.6e+02
NGC4536         |CO13-12| | 6.1e+02| 4.1e+02| 8.5e+02|
NGC4536         |NII    | | 4.1e+03| 4.0e+03| 4.3e+03|
NGC4569         |CI1-0  | | 1.4e+03| 1.2e+03| 1.6e+03|
NGC4569         |CI2-1  | | 1.2e+03| 1.1e+03| 1.2e+03|
NGC4569         |CO4-3  | | 2.0e+03| 1.8e+03| 2.2e+03|
NGC4569         |CO5-4  | | 1.5e+03| 1.4e+03| 1.7e+03|
NGC4569         |CO6-5  | | 1.0e+03| 9.8e+02| 1.1e+03|
NGC4569         |CO7-6  | | 5.7e+02| 5.2e+02| 6.2e+02|
NGC4569         |CO8-7  | | 4.5e+02| 3.9e+02| 5.0e+02|
NGC4569         |CO9-8  | | 4.1e+02| 3.1e+02| 5.2e+02|
NGC4569         |CO10-9 | | 2.5e+02| 1.6e+02| 3.3e+02|
NGC4569         |CO11-10| | 1.6e+02| 6.6e+01| 2.6e+02| 4.7e+02
NGC4569         |CO12-11| | 9.5e+01| 4.3e+01| 1.6e+02| 2.4e+02
NGC4569         |CO13-12| | 2.9e+02| 1.4e+02| 4.1e+02| 6.2e+02
NGC4569         |NII    | | 2.4e+03| 2.3e+03| 2.5e+03|
TOL1238-364     |CI1-0  | | 3.6e+02| 1.2e+02| 5.6e+02| 8.1e+02
TOL1238-364     |CI2-1  | | 2.0e+02| 1.6e+02| 2.7e+02|
TOL1238-364     |CO4-3  | | 4.3e+02| 1.4e+02| 7.4e+02| 1.2e+03
TOL1238-364     |CO5-4  | | 4.9e+02| 3.1e+02| 6.2e+02|
TOL1238-364     |CO6-5  | | 2.0e+02| 1.2e+02| 2.6e+02|
TOL1238-364     |CO7-6  | | 1.1e+02| 6.9e+01| 1.8e+02|
TOL1238-364     |CO8-7  | | 1.9e+02| 1.2e+02| 2.4e+02|
TOL1238-364     |CO9-8  | | 3.5e+02| 2.3e+02| 4.6e+02|
TOL1238-364     |CO10-9 | | 1.6e+02| 6.5e+01| 2.5e+02| 3.7e+02
TOL1238-364     |CO11-10| | 1.8e+02| 8.1e+01| 2.8e+02| 4.2e+02
TOL1238-364     |CO12-11| | 9.8e+01| 3.4e+01| 1.6e+02| 2.6e+02
TOL1238-364     |CO13-12| | 1.6e+02| 7.4e+01| 2.7e+02| 4.3e+02
TOL1238-364     |NII    | | 1.6e+03| 1.5e+03| 1.7e+03|
NGC4631         |CI1-0  | | 9.9e+02| 7.6e+02| 1.2e+03|
NGC4631         |CI2-1  | | 8.2e+02| 7.4e+02| 8.9e+02|
NGC4631         |CO4-3  | | 1.5e+03| 1.2e+03| 1.8e+03|
NGC4631         |CO5-4  | | 1.0e+03| 8.5e+02| 1.2e+03|
NGC4631         |CO6-5  | | 7.7e+02| 6.8e+02| 8.7e+02|
NGC4631         |CO7-6  | | 3.6e+02| 3.0e+02| 4.3e+02|
NGC4631         |CO9-8  | | 3.0e+02| 8.8e+01| 5.1e+02| 1.0e+03
NGC4631         |CO10-9 | | 3.8e+02| 1.4e+02| 5.7e+02| 8.3e+02
NGC4631         |CO12-11| | 2.2e+02| 6.5e+01| 3.6e+02| 5.6e+02
NGC4631         |NII    | | 1.2e+04| 1.2e+04| 1.2e+04|
NGC4710         |CI1-0  | | 1.5e+02| 4.2e+01| 2.9e+02| 4.6e+02
NGC4710         |CI2-1  | | 3.7e+02| 3.2e+02| 4.2e+02|
NGC4710         |CO4-3  | | 6.1e+02| 4.3e+02| 7.8e+02|
NGC4710         |CO5-4  | | 5.0e+02| 3.8e+02| 6.2e+02|
NGC4710         |CO6-5  | | 2.5e+02| 2.0e+02| 3.1e+02|
NGC4710         |CO7-6  | | 7.9e+01| 3.1e+01| 1.3e+02| 1.8e+02
NGC4710         |CO8-7  | | 6.0e+01| 1.2e+01| 1.0e+02| 2.2e+02
NGC4710         |CO9-8  | | 4.5e+01| 8.0e+00| 1.1e+02| 2.8e+02
NGC4710         |CO10-9 | | 9.7e+01| 3.6e+01| 1.7e+02| 3.1e+02
NGC4710         |CO11-10| | 3.3e+01| 3.9e+00| 8.2e+01| 1.8e+02
NGC4710         |CO12-11| | 1.6e+01| 3.7e-01| 5.2e+01| 1.2e+02
NGC4710         |CO13-12| | 3.5e+01| 5.6e+00| 8.8e+01| 1.9e+02
NGC4710         |NII    | | 3.5e+03| 3.4e+03| 3.6e+03|
NGC4736         |CI1-0  | | 5.9e+02| 4.9e+02| 7.0e+02|
NGC4736         |CI2-1  | | 1.1e+03| 1.0e+03| 1.1e+03|
NGC4736         |CO4-3  | | 9.1e+02| 8.0e+02| 1.0e+03|
NGC4736         |CO5-4  | | 1.1e+03| 9.7e+02| 1.2e+03|
NGC4736         |CO6-5  | | 6.1e+02| 5.6e+02| 6.8e+02|
NGC4736         |CO7-6  | | 3.7e+02| 3.2e+02| 4.2e+02|
NGC4736         |CO8-7  | | 1.2e+02| 5.3e+01| 1.9e+02| 2.8e+02
NGC4736         |CO9-8  | | 1.7e+02| 3.6e+01| 3.9e+02| 6.3e+02
NGC4736         |CO12-11| | 2.1e+02| 7.5e+01| 3.4e+02| 6.2e+02
NGC4736         |CO13-12| | 1.3e+02| 4.7e+01| 2.5e+02| 4.0e+02
NGC4736         |NII    | | 3.1e+03| 2.9e+03| 3.2e+03|
Mrk 231         |CI1-0  | | 3.8e+02| 1.6e+02| 5.8e+02| 8.4e+02
Mrk 231         |CI2-1  | | 5.1e+02| 4.5e+02| 5.5e+02|
Mrk 231         |CO5-4  | | 7.5e+02| 6.2e+02| 8.8e+02|
Mrk 231         |CO6-5  | | 9.4e+02| 8.6e+02| 1.0e+03|
Mrk 231         |CO7-6  | | 9.4e+02| 8.8e+02| 1.0e+03|
Mrk 231         |CO8-7  | | 8.2e+02| 7.7e+02| 8.8e+02|
Mrk 231         |CO9-8  | | 5.2e+02| 4.4e+02| 5.9e+02|
Mrk 231         |CO10-9 | | 7.0e+02| 6.3e+02| 7.7e+02|
Mrk 231         |CO11-10| | 5.7e+02| 5.2e+02| 6.2e+02|
Mrk 231         |CO12-11| | 4.1e+02| 3.7e+02| 4.5e+02|
Mrk 231         |CO13-12| | 3.0e+02| 2.6e+02| 3.4e+02|
Mrk 231         |NII    |X| 6.1e+02| 5.3e+02| 6.9e+02|
NGC4826         |CI1-0  | | 1.9e+03| 1.7e+03| 2.1e+03|
NGC4826         |CI2-1  | | 1.7e+03| 1.6e+03| 1.7e+03|
NGC4826         |CO4-3  | | 3.1e+03| 2.9e+03| 3.4e+03|
NGC4826         |CO5-4  | | 3.0e+03| 2.8e+03| 3.1e+03|
NGC4826         |CO6-5  | | 2.4e+03| 2.3e+03| 2.4e+03|
NGC4826         |CO7-6  | | 1.1e+03| 1.0e+03| 1.2e+03|
NGC4826         |CO8-7  | | 4.1e+02| 2.9e+02| 5.4e+02|
NGC4826         |CO9-8  | | 2.4e+02| 6.9e+01| 4.5e+02| 6.6e+02
NGC4826         |CO10-9 | | 1.6e+02| 3.4e+01| 3.0e+02| 4.9e+02
NGC4826         |CO12-11| | 6.6e+01| 7.6e-01| 1.7e+02| 3.7e+02
NGC4826         |NII    | | 8.5e+03| 8.2e+03| 8.8e+03|
MCG-02-33-098   |CI1-0  | | 3.3e+01| 4.8e+00| 9.3e+01| 1.7e+02
MCG-02-33-098   |CI2-1  | | 8.0e+01| 2.5e+01| 1.3e+02| 1.8e+02
MCG-02-33-098   |CO4-3  | | 5.7e+01| 1.7e+01| 1.5e+02| 2.0e+02
MCG-02-33-098   |CO5-4  | | 1.6e+02| 9.4e+01| 2.5e+02|
MCG-02-33-098   |CO6-5  | | 2.8e+02| 2.0e+02| 3.5e+02|
MCG-02-33-098   |CO7-6  | | 2.1e+02| 1.5e+02| 2.6e+02|
MCG-02-33-098   |CO8-7  | | 7.4e+01| 1.8e+01| 1.5e+02| 2.7e+02
MCG-02-33-098   |CO9-8  | | 1.9e+02| 6.9e+01| 3.1e+02| 4.7e+02
MCG-02-33-098   |CO10-9 | | 6.8e+01| 1.5e+01| 1.6e+02| 2.8e+02
MCG-02-33-098   |CO13-12| | 9.2e+01| 3.2e+01| 1.6e+02| 2.9e+02
MCG-02-33-098   |NII    | | 5.9e+02| 5.2e+02| 6.7e+02|
ESO507-G070     |CI1-0  | | 2.1e+02| 5.5e+01| 4.4e+02| 6.7e+02
ESO507-G070     |CI2-1  | | 5.1e+02| 4.5e+02| 5.7e+02|
ESO507-G070     |CO5-4  | | 6.5e+02| 5.5e+02| 8.0e+02|
ESO507-G070     |CO6-5  | | 7.2e+02| 6.6e+02| 7.8e+02|
ESO507-G070     |CO7-6  | | 7.3e+02| 6.7e+02| 7.9e+02|
ESO507-G070     |CO8-7  | | 7.0e+02| 6.2e+02| 7.6e+02|
ESO507-G070     |CO9-8  | | 4.7e+02| 3.9e+02| 5.4e+02|
ESO507-G070     |CO10-9 | | 3.6e+02| 2.9e+02| 4.3e+02|
ESO507-G070     |CO11-10| | 2.3e+02| 1.6e+02| 3.0e+02|
ESO507-G070     |CO12-11| | 2.0e+02| 1.5e+02| 2.5e+02|
ESO507-G070     |CO13-12| | 1.4e+02| 9.2e+01| 1.9e+02|
ESO507-G070     |NII    |X| 8.5e+02| 7.7e+02| 9.3e+02|
NGC5010         |CI1-0  | | 2.8e+02| 8.5e+01| 5.7e+02| 8.9e+02
NGC5010         |CI2-1  | | 6.9e+02| 5.9e+02| 7.7e+02|
NGC5010         |CO4-3  | | 1.6e+03| 9.9e+02| 2.1e+03|
NGC5010         |CO5-4  | | 9.1e+02| 6.1e+02| 1.2e+03|
NGC5010         |CO6-5  | | 5.8e+02| 4.4e+02| 7.0e+02|
NGC5010         |CO7-6  | | 3.4e+02| 2.4e+02| 4.4e+02|
NGC5010         |CO8-7  | | 1.8e+02| 8.1e+01| 3.0e+02| 5.0e+02
NGC5010         |CO10-9 | | 1.6e+02| 5.2e+01| 2.8e+02| 4.8e+02
NGC5010         |CO11-10| | 1.7e+02| 6.5e+01| 2.8e+02| 4.5e+02
NGC5010         |CO12-11| | 9.9e+01| 2.3e+01| 1.9e+02| 3.4e+02
NGC5010         |NII    |X| 4.6e+03| 4.4e+03| 4.8e+03|
IRAS13120-5453  |CI1-0  | | 1.4e+03| 1.2e+03| 1.8e+03|
IRAS13120-5453  |CI2-1  | | 1.7e+03| 1.6e+03| 1.8e+03|
IRAS13120-5453  |CO5-4  | | 2.4e+03| 2.2e+03| 2.6e+03|
IRAS13120-5453  |CO6-5  | | 2.3e+03| 2.2e+03| 2.4e+03|
IRAS13120-5453  |CO7-6  | | 2.1e+03| 2.0e+03| 2.2e+03|
IRAS13120-5453  |CO8-7  | | 1.8e+03| 1.6e+03| 1.9e+03|
IRAS13120-5453  |CO9-8  | | 1.1e+03| 1.0e+03| 1.2e+03|
IRAS13120-5453  |CO10-9 | | 1.1e+03| 9.7e+02| 1.2e+03|
IRAS13120-5453  |CO11-10| | 6.5e+02| 5.6e+02| 7.4e+02|
IRAS13120-5453  |CO12-11| | 4.0e+02| 3.3e+02| 4.8e+02|
IRAS13120-5453  |CO13-12| | 2.7e+02| 2.0e+02| 3.4e+02|
IRAS13120-5453  |NII    |X| 2.2e+03| 2.0e+03| 2.3e+03|
NGC5055         |CI1-0  | | 9.8e+02| 7.0e+02| 1.2e+03|
NGC5055         |CI2-1  | | 8.3e+02| 7.5e+02| 9.0e+02|
NGC5055         |CO4-3  | | 1.0e+03| 7.0e+02| 1.2e+03|
NGC5055         |CO5-4  | | 6.0e+02| 3.6e+02| 8.5e+02|
NGC5055         |CO6-5  | | 1.6e+02| 6.3e+01| 2.6e+02| 4.4e+02
NGC5055         |CO7-6  | | 1.2e+02| 4.8e+01| 2.1e+02| 3.1e+02
NGC5055         |CO8-7  | | 2.0e+02| 1.1e+02| 3.0e+02| 4.3e+02
NGC5055         |CO9-8  | | 1.0e+02| 7.8e+00| 2.5e+02| 4.9e+02
NGC5055         |CO11-10| | 2.3e+02| 6.8e+01| 4.2e+02| 7.5e+02
NGC5055         |CO12-11| | 7.2e+01| 6.0e+00| 1.7e+02| 2.9e+02
NGC5055         |NII    | | 6.7e+03| 6.4e+03| 7.0e+03|
Arp193          |CI1-0  | | 1.1e+03| 8.1e+02| 1.4e+03|
Arp193          |CI2-1  | | 1.1e+03| 1.0e+03| 1.1e+03|
Arp193          |CO5-4  | | 1.8e+03| 1.7e+03| 1.9e+03|
Arp193          |CO6-5  | | 1.6e+03| 1.5e+03| 1.6e+03|
Arp193          |CO7-6  | | 9.9e+02| 9.5e+02| 1.0e+03|
Arp193          |CO8-7  | | 6.4e+02| 6.0e+02| 6.8e+02|
Arp193          |CO9-8  | | 4.8e+02| 4.4e+02| 5.3e+02|
Arp193          |CO10-9 | | 3.8e+02| 3.4e+02| 4.1e+02|
Arp193          |CO11-10| | 2.5e+02| 2.2e+02| 2.8e+02|
Arp193          |CO12-11| | 1.3e+02| 1.0e+02| 1.6e+02|
Arp193          |CO13-12| | 8.9e+01| 5.9e+01| 1.1e+02|
Arp193          |NII    |X| 1.4e+03| 1.4e+03| 1.5e+03|
NGC5104         |CI1-0  | | 9.4e+01| 1.5e+01| 2.5e+02| 4.6e+02
NGC5104         |CI2-1  | | 5.0e+02| 4.4e+02| 5.6e+02|
NGC5104         |CO5-4  | | 5.0e+02| 3.4e+02| 6.4e+02|
NGC5104         |CO6-5  | | 4.4e+02| 3.7e+02| 5.1e+02|
NGC5104         |CO7-6  | | 2.6e+02| 2.0e+02| 3.2e+02|
NGC5104         |CO8-7  | | 1.3e+02| 3.7e+01| 2.2e+02| 3.4e+02
NGC5104         |CO9-8  | | 1.5e+02| 4.7e+01| 2.6e+02| 4.2e+02
NGC5104         |CO10-9 | | 8.6e+01| 2.2e+01| 1.5e+02| 2.6e+02
NGC5104         |CO11-10| | 1.4e+02| 6.7e+01| 2.2e+02| 3.5e+02
NGC5104         |CO12-11| | 7.0e+01| 2.0e+01| 1.3e+02| 2.4e+02
NGC5104         |NII    |X| 1.6e+03| 1.5e+03| 1.7e+03|
MCG-03-34-064   |CI2-1  | | 1.3e+02| 6.6e+01| 1.9e+02|
MCG-03-34-064   |CO4-3  | | 3.1e+01| 5.7e+00| 6.6e+01| 1.5e+02
MCG-03-34-064   |CO5-4  | | 6.7e+01| 1.7e+01| 1.3e+02| 2.5e+02
MCG-03-34-064   |CO6-5  | | 1.4e+02| 9.3e+01| 1.9e+02|
MCG-03-34-064   |CO7-6  | | 1.4e+02| 7.0e+01| 2.0e+02|
MCG-03-34-064   |CO8-7  | | 9.2e+01| 2.6e+01| 1.6e+02| 2.7e+02
MCG-03-34-064   |CO10-9 | | 3.3e+02| 2.5e+02| 4.1e+02|
MCG-03-34-064   |CO11-10| | 1.6e+02| 9.3e+01| 2.2e+02|
MCG-03-34-064   |CO12-11| | 1.6e+02| 7.2e+01| 2.2e+02|
MCG-03-34-064   |CO13-12| | 1.6e+02| 9.6e+01| 2.3e+02|
MCG-03-34-064   |NII    |X| 4.5e+02| 3.6e+02| 5.4e+02|
Cen A           |CI1-0  | | 4.0e+03| 3.8e+03| 4.2e+03|
Cen A           |CI2-1  | | 9.5e+03| 9.3e+03| 9.6e+03|
Cen A           |CO4-3  | | 4.2e+03| 4.0e+03| 4.5e+03|
Cen A           |CO5-4  | | 3.9e+03| 3.7e+03| 4.1e+03|
Cen A           |CO6-5  | | 2.6e+03| 2.5e+03| 2.7e+03|
Cen A           |CO7-6  | | 1.6e+03| 1.4e+03| 1.7e+03|
Cen A           |CO8-7  | | 1.3e+03| 1.0e+03| 1.5e+03|
Cen A           |CO9-8  | | 9.0e+02| 3.7e+02| 1.2e+03| 1.7e+03
Cen A           |CO10-9 | | 4.8e+02| 2.8e+02| 6.8e+02| 9.7e+02
Cen A           |CO11-10| | 1.4e+02| 8.3e+00| 3.7e+02| 7.4e+02
Cen A           |CO12-11| | 2.9e+02| 1.0e+02| 4.9e+02| 7.6e+02
Cen A           |CO13-12| | 4.9e+02| 1.7e+02| 9.4e+02| 1.7e+03
Cen A           |NII    | | 1.1e+04| 1.0e+04| 1.1e+04|
NGC5135         |CI1-0  | | 1.8e+03| 1.6e+03| 2.0e+03|
NGC5135         |CI2-1  | | 1.9e+03| 1.9e+03| 1.9e+03|
NGC5135         |CO4-3  | | 2.1e+03| 1.8e+03| 2.3e+03|
NGC5135         |CO5-4  | | 1.8e+03| 1.7e+03| 1.9e+03|
NGC5135         |CO6-5  | | 1.5e+03| 1.5e+03| 1.6e+03|
NGC5135         |CO7-6  | | 9.3e+02| 8.9e+02| 9.7e+02|
NGC5135         |CO8-7  | | 6.0e+02| 5.5e+02| 6.5e+02|
NGC5135         |CO9-8  | | 4.4e+02| 3.8e+02| 5.0e+02|
NGC5135         |CO10-9 | | 3.1e+02| 2.6e+02| 3.6e+02|
NGC5135         |CO11-10| | 1.7e+02| 1.3e+02| 2.1e+02|
NGC5135         |CO12-11| | 1.7e+02| 1.4e+02| 2.0e+02|
NGC5135         |NII    | | 3.2e+03| 3.1e+03| 3.2e+03|
ESO 173-G015    |CI1-0  | | 1.6e+03| 1.3e+03| 1.8e+03|
ESO 173-G015    |CI2-1  | | 3.0e+03| 3.0e+03| 3.1e+03|
ESO 173-G015    |CO4-3  | | 4.0e+03| 3.6e+03| 4.4e+03|
ESO 173-G015    |CO5-4  | | 4.8e+03| 4.6e+03| 5.0e+03|
ESO 173-G015    |CO6-5  | | 4.8e+03| 4.7e+03| 4.9e+03|
ESO 173-G015    |CO7-6  | | 3.7e+03| 3.6e+03| 3.8e+03|
ESO 173-G015    |CO8-7  | | 3.2e+03| 3.0e+03| 3.3e+03|
ESO 173-G015    |CO9-8  | | 3.1e+03| 2.9e+03| 3.3e+03|
ESO 173-G015    |CO10-9 | | 2.6e+03| 2.5e+03| 2.8e+03|
ESO 173-G015    |CO11-10| | 2.2e+03| 2.0e+03| 2.3e+03|
ESO 173-G015    |CO12-11| | 1.4e+03| 1.3e+03| 1.5e+03|
ESO 173-G015    |CO13-12| | 9.9e+02| 8.4e+02| 1.1e+03|
ESO 173-G015    |NII    | | 3.2e+03| 3.0e+03| 3.3e+03|
NGC5194         |CI1-0  | | 1.5e+03| 1.2e+03| 1.8e+03|
NGC5194         |CI2-1  | | 2.8e+03| 2.7e+03| 2.9e+03|
NGC5194         |CO4-3  | | 1.6e+03| 1.3e+03| 1.8e+03|
NGC5194         |CO5-4  | | 1.9e+03| 1.6e+03| 2.2e+03|
NGC5194         |CO6-5  | | 1.3e+03| 1.2e+03| 1.5e+03|
NGC5194         |CO7-6  | | 8.8e+02| 7.8e+02| 9.9e+02|
NGC5194         |CO8-7  | | 4.0e+02| 2.2e+02| 5.7e+02| 7.3e+02
NGC5194         |CO9-8  | | 6.6e+02| 1.8e+02| 1.1e+03| 1.8e+03
NGC5194         |CO10-9 | | 9.0e+02| 6.3e+02| 1.2e+03| 1.8e+03
NGC5194         |CO11-10| | 5.9e+02| 2.9e+02| 8.8e+02| 1.2e+03
NGC5194         |CO12-11| | 3.1e+02| 7.8e+01| 5.7e+02| 1.0e+03
NGC5194         |CO13-12| | 5.6e+02| 1.6e+02| 1.0e+03| 1.9e+03
NGC5194         |NII    | | 2.6e+04| 2.5e+04| 2.6e+04|
IC4280          |CI1-0  | | 2.3e+02| 6.9e+01| 4.1e+02| 7.3e+02
IC4280          |CI2-1  | | 3.8e+02| 3.0e+02| 4.4e+02|
IC4280          |CO4-3  | | 7.9e+02| 5.4e+02| 1.0e+03|
IC4280          |CO5-4  | | 5.4e+02| 3.9e+02| 7.1e+02|
IC4280          |CO6-5  | | 3.5e+02| 2.6e+02| 4.2e+02|
IC4280          |CO7-6  | | 1.5e+02| 7.3e+01| 2.2e+02|
IC4280          |CO8-7  | | 1.9e+02| 9.7e+01| 2.7e+02| 4.0e+02
IC4280          |CO10-9 | | 1.9e+02| 9.8e+01| 3.0e+02| 4.6e+02
IC4280          |CO13-12| | 4.8e+01| 9.2e+00| 1.1e+02| 2.2e+02
IC4280          |NII    | | 3.4e+03| 3.2e+03| 3.4e+03|
M83             |CI1-0  | | 3.5e+03| 3.1e+03| 3.9e+03|
M83             |CI2-1  | | 4.6e+03| 4.4e+03| 4.7e+03|
M83             |CO4-3  | | 8.5e+03| 8.0e+03| 9.0e+03|
M83             |CO5-4  | | 9.5e+03| 9.1e+03| 9.9e+03|
M83             |CO6-5  | | 7.3e+03| 7.0e+03| 7.5e+03|
M83             |CO7-6  | | 4.5e+03| 4.3e+03| 4.6e+03|
M83             |CO8-7  | | 3.0e+03| 2.8e+03| 3.2e+03|
M83             |CO9-8  | | 1.5e+03| 6.7e+02| 2.0e+03| 2.7e+03
M83             |CO10-9 | | 1.2e+03| 8.4e+02| 1.5e+03|
M83             |CO11-10| | 8.5e+02| 5.5e+02| 1.2e+03|
M83             |CO12-11| | 4.3e+02| 7.0e+01| 7.7e+02| 1.3e+03
M83             |NII    | | 1.9e+04| 1.8e+04| 2.0e+04|
Mrk 273         |CI1-0  | | 3.7e+02| 1.1e+02| 5.8e+02| 1.1e+03
Mrk 273         |CI2-1  | | 6.4e+02| 5.8e+02| 6.9e+02|
Mrk 273         |CO5-4  | | 1.2e+03| 1.0e+03| 1.4e+03|
Mrk 273         |CO6-5  | | 1.2e+03| 1.1e+03| 1.3e+03|
Mrk 273         |CO7-6  | | 1.1e+03| 1.0e+03| 1.1e+03|
Mrk 273         |CO8-7  | | 7.4e+02| 6.8e+02| 7.9e+02|
Mrk 273         |CO9-8  |X| 9.4e+02| 8.3e+02| 1.0e+03|
Mrk 273         |CO10-9 |X| 1.1e+03| 1.1e+03| 1.2e+03|
Mrk 273         |CO11-10|X| 5.6e+02| 4.7e+02| 6.4e+02|
Mrk 273         |CO12-11|X| 5.1e+02| 4.2e+02| 5.9e+02|
Mrk 273         |CO13-12|X| 5.7e+02| 4.9e+02| 6.6e+02|
Mrk 273         |NII    |X| 1.0e+03| 9.5e+02| 1.1e+03|
4C 12.50        |CI2-1  | | 4.0e+01| 9.0e+00| 8.4e+01| 1.7e+02
4C 12.50        |CO5-4  | | 2.3e+02| 9.2e+01| 4.0e+02| 6.1e+02
4C 12.50        |CO6-5  | | 1.0e+02| 2.7e+01| 2.1e+02| 3.5e+02
4C 12.50        |CO7-6  | | 9.0e+01| 3.9e+01| 1.5e+02|
4C 12.50        |CO8-7  | | 4.7e+01| 1.6e+01| 9.6e+01| 1.6e+02
4C 12.50        |CO10-9 | | 7.9e+01| 3.0e+01| 1.3e+02| 2.2e+02
4C 12.50        |CO11-10| | 5.0e+01| 1.5e+01| 9.5e+01| 1.7e+02
4C 12.50        |CO12-11| | 4.0e+01| 1.0e+01| 8.2e+01| 1.3e+02
4C 12.50        |CO13-12| | 2.7e+01| 6.7e+00| 6.8e+01| 1.1e+02
4C 12.50        |NII    | | 3.6e+01| 7.7e+00| 7.8e+01| 1.3e+02
UGC08739        |CI1-0  | | 3.6e+02| 1.2e+02| 5.2e+02| 7.8e+02
UGC08739        |CI2-1  | | 4.8e+02| 4.3e+02| 5.4e+02|
UGC08739        |CO4-3  | | 3.3e+02| 8.4e+01| 4.9e+02| 7.1e+02
UGC08739        |CO5-4  | | 6.2e+02| 4.9e+02| 7.5e+02|
UGC08739        |CO6-5  | | 2.2e+02| 1.4e+02| 2.9e+02|
UGC08739        |CO7-6  | | 1.8e+02| 1.3e+02| 2.5e+02|
UGC08739        |CO8-7  | | 2.8e+02| 2.0e+02| 3.6e+02|
UGC08739        |CO9-8  | | 2.3e+02| 1.0e+02| 3.4e+02| 5.3e+02
UGC08739        |CO10-9 | | 9.5e+01| 2.6e+01| 2.0e+02| 3.5e+02
UGC08739        |CO11-10| | 1.4e+02| 4.7e+01| 2.5e+02| 4.3e+02
UGC08739        |CO13-12| | 7.5e+01| 1.3e+01| 1.7e+02| 2.9e+02
UGC08739        |NII    | | 2.0e+03| 2.0e+03| 2.1e+03|
ESO221-IG010    |CI1-0  | | 2.1e+02| 5.9e+01| 3.5e+02| 5.9e+02
ESO221-IG010    |CI2-1  | | 3.3e+02| 2.4e+02| 4.1e+02|
ESO221-IG010    |CO4-3  | | 8.3e+01| 1.0e+01| 2.6e+02| 4.8e+02
ESO221-IG010    |CO5-4  | | 5.7e+02| 4.6e+02| 6.9e+02|
ESO221-IG010    |CO6-5  | | 4.1e+02| 3.3e+02| 4.9e+02|
ESO221-IG010    |CO7-6  | | 2.6e+02| 1.8e+02| 3.5e+02|
ESO221-IG010    |CO8-7  | | 9.8e+01| 2.0e+01| 2.1e+02| 5.3e+02
ESO221-IG010    |CO9-8  | | 3.2e+02| 1.6e+02| 4.9e+02| 8.4e+02
ESO221-IG010    |CO10-9 | | 1.8e+02| 5.0e+01| 3.2e+02| 5.4e+02
ESO221-IG010    |CO13-12| | 2.2e+02| 9.4e+01| 3.6e+02| 5.5e+02
ESO221-IG010    |NII    | | 3.3e+03| 3.2e+03| 3.5e+03|
Mrk 463         |CI1-0  | | 1.4e+02| 3.4e+01| 2.9e+02| 5.0e+02
Mrk 463         |CI2-1  | | 1.1e+02| 6.9e+01| 1.5e+02|
Mrk 463         |CO5-4  | | 9.6e+01| 2.2e+01| 2.1e+02| 3.7e+02
Mrk 463         |CO6-5  | | 1.9e+02| 1.4e+02| 2.5e+02|
Mrk 463         |CO7-6  | | 1.1e+02| 7.0e+01| 1.4e+02|
Mrk 463         |CO8-7  | | 8.8e+01| 4.1e+01| 1.3e+02| 2.0e+02
Mrk 463         |CO9-8  | | 4.5e+01| 1.0e+01| 1.1e+02| 1.9e+02
Mrk 463         |CO10-9 | | 3.7e+01| 7.4e+00| 7.8e+01| 1.2e+02
Mrk 463         |CO11-10| | 6.6e+01| 2.6e+01| 1.2e+02| 1.7e+02
Mrk 463         |CO12-11| | 5.0e+01| 1.8e+01| 1.0e+02| 1.6e+02
Mrk 463         |NII    | | 1.0e+02| 6.4e+01| 1.6e+02|
M101_02         |CI1-0  | | 1.7e+02| 4.4e+01| 3.2e+02| 5.2e+02
M101_02         |CI2-1  | | 1.1e+02| 3.1e+01| 1.8e+02| 2.8e+02
M101_02         |CO4-3  | | 5.4e+02| 2.8e+02| 8.2e+02| 1.1e+03
M101_02         |CO5-4  | | 1.6e+02| 3.2e+01| 3.0e+02| 5.8e+02
M101_02         |CO6-5  | | 7.8e+01| 2.8e+01| 1.8e+02| 2.7e+02
M101_02         |CO7-6  | | 1.8e+02| 8.8e+01| 2.5e+02|
M101_02         |CO8-7  | | 6.5e+01| 1.6e+01| 1.3e+02| 2.8e+02
M101_02         |CO9-8  | | 2.2e+02| 1.0e+02| 3.5e+02| 5.3e+02
M101_02         |CO10-9 | | 9.7e+01| 1.6e+01| 2.0e+02| 3.3e+02
M101_02         |CO11-10| | 1.3e+02| 3.8e+01| 2.7e+02| 4.0e+02
M101_02         |CO12-11| | 8.4e+01| 2.6e+01| 1.6e+02| 2.7e+02
M101_02         |NII    | | 1.7e+03| 1.6e+03| 1.8e+03|
OQ 208          |CI1-0  | | 5.3e+02| 3.2e+02| 7.4e+02|
OQ 208          |CI2-1  | | 5.9e+01| 2.8e+01| 9.8e+01| 1.6e+02
OQ 208          |CO5-4  | | 2.6e+02| 1.5e+02| 4.2e+02| 6.4e+02
OQ 208          |CO7-6  | | 5.0e+01| 2.0e+01| 9.2e+01| 1.4e+02
OQ 208          |CO8-7  | | 4.7e+01| 1.4e+01| 9.1e+01| 1.5e+02
OQ 208          |CO10-9 | | 2.5e+02| 6.9e+01| 4.8e+02| 7.7e+02
OQ 208          |CO12-11| | 4.8e+02| 2.7e+02| 6.8e+02|
OQ 208          |CO13-12| | 1.2e+02| 2.1e+01| 2.2e+02| 3.5e+02
OQ 208          |NII    | | 4.2e+02| 2.7e+02| 5.7e+02|
NGC5653         |CI1-0  | | 3.2e+02| 5.9e+01| 6.0e+02| 8.6e+02
NGC5653         |CI2-1  | | 5.3e+02| 4.0e+02| 6.5e+02|
NGC5653         |CO4-3  | | 5.6e+02| 1.9e+02| 8.7e+02| 1.2e+03
NGC5653         |CO5-4  | | 1.2e+03| 1.1e+03| 1.4e+03|
NGC5653         |CO6-5  | | 4.9e+02| 3.5e+02| 6.3e+02|
NGC5653         |CO7-6  | | 1.6e+02| 5.5e+01| 2.7e+02| 3.8e+02
NGC5653         |CO8-7  | | 3.6e+02| 2.2e+02| 5.2e+02|
NGC5653         |CO9-8  | | 1.5e+02| 3.5e+01| 3.0e+02| 5.6e+02
NGC5653         |CO10-9 | | 7.9e+01| 1.1e+01| 2.0e+02| 3.5e+02
NGC5653         |CO11-10| | 1.3e+02| 1.8e+01| 2.6e+02| 4.8e+02
NGC5653         |CO12-11| | 5.6e+01| 6.3e+00| 1.4e+02| 3.0e+02
NGC5653         |CO13-12| | 1.2e+02| 2.8e+01| 2.8e+02| 5.1e+02
NGC5653         |NII    | | 4.7e+03| 4.5e+03| 4.9e+03|
IRAS 14348-1447 |CI2-1  | | 3.6e+02| 3.0e+02| 4.1e+02|
IRAS 14348-1447 |CO5-4  | | 3.1e+02| 1.4e+02| 5.2e+02| 7.8e+02
IRAS 14348-1447 |CO6-5  | | 3.4e+02| 2.4e+02| 4.2e+02|
IRAS 14348-1447 |CO7-6  | | 3.1e+02| 2.6e+02| 3.6e+02|
IRAS 14348-1447 |CO8-7  | | 4.3e+02| 3.7e+02| 4.9e+02|
IRAS 14348-1447 |CO9-8  | | 1.3e+02| 6.7e+01| 1.9e+02| 3.0e+02
IRAS 14348-1447 |CO10-9 | | 2.6e+02| 2.0e+02| 3.2e+02|
IRAS 14348-1447 |CO11-10| | 1.7e+02| 1.2e+02| 2.2e+02|
IRAS 14348-1447 |CO12-11| | 5.6e+01| 1.6e+01| 1.0e+02| 1.7e+02
IRAS 14348-1447 |CO13-12| | 1.5e+02| 1.2e+02| 1.9e+02|
IRAS 14348-1447 |NII    | | 2.4e+02| 2.1e+02| 2.8e+02|
NGC5713         |CI1-0  | | 6.7e+02| 5.1e+02| 8.3e+02|
NGC5713         |CI2-1  | | 6.6e+02| 6.0e+02| 7.2e+02|
NGC5713         |CO4-3  | | 1.3e+03| 1.2e+03| 1.5e+03|
NGC5713         |CO5-4  | | 1.3e+03| 1.1e+03| 1.4e+03|
NGC5713         |CO6-5  | | 9.4e+02| 8.6e+02| 1.0e+03|
NGC5713         |CO7-6  | | 5.9e+02| 5.3e+02| 6.5e+02|
NGC5713         |CO8-7  | | 2.8e+02| 2.0e+02| 3.4e+02|
NGC5713         |CO9-8  | | 1.8e+02| 7.5e+01| 3.1e+02| 5.6e+02
NGC5713         |CO10-9 | | 1.6e+02| 5.0e+01| 2.8e+02| 4.6e+02
NGC5713         |CO11-10| | 3.1e+02| 1.6e+02| 4.4e+02| 6.7e+02
NGC5713         |CO12-11| | 6.6e+01| 9.9e+00| 1.5e+02| 2.7e+02
NGC5713         |CO13-12| | 2.7e+02| 8.3e+01| 4.5e+02| 6.6e+02
NGC5713         |NII    | | 4.7e+03| 4.5e+03| 4.9e+03|
IRAS 14378-3651 |CI1-0  | | 1.0e+03| 7.4e+02| 1.2e+03|
IRAS 14378-3651 |CI2-1  | | 1.7e+02| 1.3e+02| 2.3e+02|
IRAS 14378-3651 |CO5-4  | | 4.2e+02| 2.4e+02| 6.1e+02|
IRAS 14378-3651 |CO6-5  | | 2.7e+02| 1.9e+02| 3.7e+02|
IRAS 14378-3651 |CO7-6  | | 4.1e+02| 3.6e+02| 4.6e+02|
IRAS 14378-3651 |CO8-7  | | 2.3e+02| 1.8e+02| 2.9e+02|
IRAS 14378-3651 |CO9-8  | | 1.9e+02| 9.7e+01| 3.0e+02| 4.6e+02
IRAS 14378-3651 |CO10-9 | | 1.2e+02| 6.8e+01| 2.0e+02|
IRAS 14378-3651 |CO11-10| | 1.4e+02| 7.2e+01| 2.0e+02|
IRAS 14378-3651 |CO12-11| | 1.3e+02| 8.1e+01| 1.8e+02|
IRAS 14378-3651 |CO13-12| | 1.1e+02| 5.6e+01| 1.5e+02|
Mrk 478         |CI1-0  | | 3.1e+02| 1.0e+02| 5.2e+02| 6.7e+02
Mrk 478         |CI2-1  | | 8.6e+01| 4.4e+01| 1.4e+02| 2.0e+02
Mrk 478         |CO6-5  | | 8.6e+01| 2.3e+01| 2.0e+02| 2.9e+02
Mrk 478         |CO7-6  | | 4.2e+01| 7.7e+00| 9.2e+01| 1.5e+02
Mrk 478         |CO9-8  | | 4.5e+01| 9.4e+00| 8.9e+01| 1.4e+02
Mrk 478         |CO11-10| | 6.7e+01| 3.2e+01| 1.1e+02| 1.6e+02
Mrk 478         |CO12-11| | 4.6e+01| 1.2e+01| 8.9e+01| 1.6e+02
Mrk 478         |CO13-12| | 4.1e+01| 8.4e+00| 7.4e+01| 1.1e+02
Mrk 478         |NII    | | 3.2e+01| 6.5e+00| 7.8e+01| 1.4e+02
NGC5734a        |CI1-0  | | 2.8e+02| 8.2e+01| 4.8e+02| 9.1e+02
NGC5734a        |CI2-1  | | 4.9e+02| 3.9e+02| 5.9e+02|
NGC5734a        |CO4-3  | | 4.6e+02| 2.6e+02| 7.4e+02|
NGC5734a        |CO5-4  | | 4.3e+02| 2.2e+02| 7.0e+02| 1.1e+03
NGC5734a        |CO6-5  | | 2.2e+02| 9.3e+01| 3.3e+02| 5.0e+02
NGC5734a        |CO7-6  | | 1.1e+02| 3.4e+01| 2.2e+02| 3.2e+02
NGC5734a        |CO8-7  | | 2.7e+02| 1.6e+02| 3.9e+02| 7.0e+02
NGC5734a        |CO9-8  | | 1.3e+02| 3.7e+01| 2.4e+02| 4.5e+02
NGC5734a        |CO10-9 | | 1.3e+02| 4.0e+01| 2.6e+02| 4.8e+02
NGC5734a        |CO11-10| | 1.8e+02| 6.3e+01| 3.1e+02| 5.2e+02
NGC5734a        |CO12-11| | 1.6e+02| 7.2e+01| 2.7e+02| 4.7e+02
NGC5734a        |CO13-12| | 9.6e+01| 1.9e+01| 2.2e+02| 4.3e+02
NGC5734a        |NII    | | 3.7e+03| 3.6e+03| 3.9e+03|
3C 305          |CO9-8  | | 1.0e+02| 2.9e+01| 2.0e+02| 3.7e+02
3C 305          |CO10-9 | | 1.4e+02| 4.1e+01| 2.6e+02| 4.3e+02
3C 305          |CO11-10| | 1.3e+02| 3.7e+01| 2.3e+02| 3.7e+02
3C 305          |CO12-11| | 1.4e+02| 4.0e+01| 2.2e+02| 4.0e+02
3C 305          |NII    | | 3.5e+02| 2.5e+02| 4.6e+02|
VV340a          |CI1-0  | | 1.1e+03| 8.6e+02| 1.3e+03|
VV340a          |CI2-1  | | 6.3e+02| 5.8e+02| 6.9e+02|
VV340a          |CO5-4  | | 4.9e+02| 3.4e+02| 6.8e+02|
VV340a          |CO6-5  | | 4.1e+02| 3.3e+02| 5.0e+02|
VV340a          |CO7-6  | | 1.8e+02| 1.3e+02| 2.3e+02|
VV340a          |CO8-7  | | 1.1e+02| 4.1e+01| 1.8e+02| 2.9e+02
VV340a          |CO9-8  | | 7.8e+01| 1.9e+01| 1.5e+02| 3.0e+02
VV340a          |CO10-9 | | 9.1e+01| 3.7e+01| 1.5e+02| 2.8e+02
VV340a          |CO11-10| | 5.1e+01| 8.2e+00| 1.0e+02| 1.6e+02
VV340a          |CO13-12| | 6.4e+01| 2.0e+01| 1.2e+02| 2.1e+02
VV340a          |NII    |X| 3.8e+03| 3.7e+03| 3.9e+03|
IC4518ABa       |CI1-0  | | 1.4e+02| 6.4e+01| 2.4e+02| 3.5e+02
IC4518ABa       |CI2-1  | | 5.2e+02| 4.6e+02| 5.8e+02|
IC4518ABa       |CO4-3  | | 2.2e+02| 7.5e+01| 3.8e+02| 6.0e+02
IC4518ABa       |CO5-4  | | 3.8e+02| 3.0e+02| 4.7e+02|
IC4518ABa       |CO6-5  | | 3.1e+02| 2.5e+02| 3.8e+02|
IC4518ABa       |CO7-6  | | 1.7e+02| 1.2e+02| 2.2e+02|
IC4518ABa       |CO8-7  | | 1.9e+02| 1.3e+02| 2.7e+02|
IC4518ABa       |CO9-8  | | 2.1e+02| 8.1e+01| 3.2e+02| 4.6e+02
IC4518ABa       |CO10-9 | | 6.3e+01| 1.7e+01| 1.3e+02| 2.6e+02
IC4518ABa       |CO11-10| | 2.7e+02| 1.9e+02| 3.6e+02|
IC4518ABa       |NII    | | 6.9e+02| 6.1e+02| 7.8e+02|
NGC5866         |CI1-0  | | 3.2e+02| 9.1e+01| 5.3e+02| 8.0e+02
NGC5866         |CI2-1  | | 4.5e+02| 4.0e+02| 5.0e+02|
NGC5866         |CO4-3  | | 8.5e+02| 5.5e+02| 1.2e+03|
NGC5866         |CO5-4  | | 4.5e+02| 3.3e+02| 6.2e+02|
NGC5866         |CO6-5  | | 3.2e+02| 2.4e+02| 4.0e+02|
NGC5866         |CO7-6  | | 1.8e+02| 1.2e+02| 2.4e+02|
NGC5866         |CO8-7  | | 2.7e+02| 1.8e+02| 3.7e+02|
NGC5866         |CO9-8  | | 5.8e+01| 1.3e+01| 1.1e+02| 2.4e+02
NGC5866         |CO10-9 | | 6.1e+01| 1.4e+01| 1.2e+02| 2.3e+02
NGC5866         |CO11-10| | 4.8e+01| 1.1e+01| 1.0e+02| 2.3e+02
NGC5866         |NII    | | 1.2e+03| 1.2e+03| 1.3e+03|
CGCG049-057     |CI1-0  | | 5.3e+02| 3.1e+02| 7.4e+02| 1.1e+03
CGCG049-057     |CI2-1  | | 4.3e+02| 3.6e+02| 4.8e+02|
CGCG049-057     |CO4-3  | | 7.6e+02| 5.2e+02| 9.6e+02|
CGCG049-057     |CO5-4  | | 8.6e+02| 7.3e+02| 9.7e+02|
CGCG049-057     |CO6-5  | | 1.0e+03| 9.5e+02| 1.1e+03|
CGCG049-057     |CO7-6  | | 9.7e+02| 9.1e+02| 1.0e+03|
CGCG049-057     |CO8-7  | | 7.1e+02| 6.2e+02| 7.7e+02|
CGCG049-057     |CO9-8  | | 5.8e+02| 5.0e+02| 6.7e+02|
CGCG049-057     |CO10-9 | | 6.3e+02| 5.5e+02| 7.2e+02|
CGCG049-057     |CO11-10| | 2.7e+02| 2.2e+02| 3.1e+02|
CGCG049-057     |CO12-11| | 1.3e+02| 8.1e+01| 1.7e+02|
CGCG049-057     |CO13-12| | 7.0e+01| 2.6e+01| 1.2e+02| 2.4e+02
CGCG049-057     |NII    | | 4.5e+02| 4.0e+02| 5.1e+02|
3C 315          |CO10-9 | | 4.8e+01| 1.3e+01| 8.9e+01| 1.4e+02
3C 315          |CO11-10| | 4.3e+01| 1.2e+01| 8.5e+01| 1.4e+02
3C 315          |CO12-11| | 4.4e+01| 1.1e+01| 8.4e+01| 1.4e+02
3C 315          |NII    | | 7.5e+01| 3.5e+01| 1.1e+02| 1.6e+02
VV705           |CI1-0  | | 3.2e+02| 1.3e+02| 6.3e+02| 1.0e+03
VV705           |CI2-1  | | 3.2e+02| 2.7e+02| 3.8e+02|
VV705           |CO5-4  | | 5.6e+02| 3.8e+02| 7.3e+02|
VV705           |CO6-5  | | 3.0e+02| 2.1e+02| 3.9e+02|
VV705           |CO7-6  | | 3.5e+02| 3.0e+02| 4.0e+02|
VV705           |CO8-7  | | 2.5e+02| 1.9e+02| 3.2e+02|
VV705           |CO9-8  | | 1.6e+02| 8.9e+01| 2.4e+02| 3.6e+02
VV705           |CO10-9 | | 1.4e+02| 7.8e+01| 2.0e+02|
VV705           |CO11-10| | 1.3e+02| 8.7e+01| 1.7e+02|
VV705           |CO12-11| | 1.3e+02| 8.3e+01| 1.8e+02|
VV705           |CO13-12| | 9.9e+01| 5.5e+01| 1.5e+02|
VV705           |NII    | | 4.6e+02| 4.1e+02| 5.0e+02|
ESO099-G004     |CI1-0  | | 2.5e+02| 6.5e+01| 4.5e+02| 9.5e+02
ESO099-G004     |CI2-1  | | 3.3e+02| 3.0e+02| 3.7e+02|
ESO099-G004     |CO5-4  | | 4.5e+02| 2.8e+02| 6.1e+02|
ESO099-G004     |CO6-5  | | 4.9e+02| 4.3e+02| 5.6e+02|
ESO099-G004     |CO7-6  | | 3.3e+02| 2.9e+02| 3.7e+02|
ESO099-G004     |CO8-7  | | 1.4e+02| 9.8e+01| 1.8e+02|
ESO099-G004     |CO9-8  | | 3.5e+02| 2.9e+02| 4.2e+02|
ESO099-G004     |CO10-9 | | 1.7e+02| 1.1e+02| 2.3e+02|
ESO099-G004     |CO11-10| | 1.4e+02| 9.5e+01| 2.0e+02|
ESO099-G004     |CO12-11| | 8.9e+01| 5.0e+01| 1.3e+02| 1.9e+02
ESO099-G004     |CO13-12| | 1.4e+02| 8.8e+01| 1.9e+02|
ESO099-G004     |NII    |X| 1.7e+03| 1.6e+03| 1.7e+03|
IRAS 15250+3609 |CI1-0  | | 4.7e+02| 2.4e+02| 7.7e+02| 1.1e+03
IRAS 15250+3609 |CI2-1  | | 1.0e+02| 5.0e+01| 1.6e+02| 2.6e+02
IRAS 15250+3609 |CO5-4  | | 1.9e+02| 5.0e+01| 3.6e+02| 5.2e+02
IRAS 15250+3609 |CO6-5  | | 2.8e+02| 1.9e+02| 3.8e+02|
IRAS 15250+3609 |CO7-6  | | 2.8e+02| 2.2e+02| 3.3e+02|
IRAS 15250+3609 |CO8-7  | | 2.1e+02| 1.3e+02| 2.7e+02| 3.6e+02
IRAS 15250+3609 |CO9-8  | | 9.3e+01| 2.9e+01| 1.7e+02| 3.0e+02
IRAS 15250+3609 |CO10-9 | | 1.4e+02| 7.5e+01| 2.0e+02| 2.9e+02
IRAS 15250+3609 |CO11-10| | 1.1e+02| 4.2e+01| 1.6e+02| 2.5e+02
IRAS 15250+3609 |CO12-11| | 9.3e+01| 4.2e+01| 1.6e+02| 2.3e+02
IRAS 15250+3609 |NII    | | 8.8e+01| 3.4e+01| 1.4e+02| 2.1e+02
NGC5936         |CI1-0  | | 2.5e+02| 7.0e+01| 4.3e+02| 7.5e+02
NGC5936         |CI2-1  | | 4.4e+02| 3.6e+02| 5.2e+02|
NGC5936         |CO4-3  | | 3.8e+02| 1.6e+02| 5.8e+02| 9.5e+02
NGC5936         |CO5-4  | | 6.1e+02| 4.3e+02| 7.8e+02|
NGC5936         |CO6-5  | | 5.3e+02| 4.4e+02| 6.3e+02|
NGC5936         |CO7-6  | | 2.5e+02| 1.5e+02| 3.3e+02|
NGC5936         |CO8-7  | | 3.7e+02| 2.4e+02| 4.8e+02|
NGC5936         |CO9-8  | | 3.3e+02| 1.4e+02| 5.4e+02| 8.6e+02
NGC5936         |CO10-9 | | 1.6e+02| 5.1e+01| 3.1e+02| 5.7e+02
NGC5936         |CO12-11| | 2.1e+02| 6.4e+01| 3.9e+02| 6.3e+02
NGC5936         |NII    | | 2.5e+03| 2.3e+03| 2.6e+03|
Arp220          |CI1-0  | | 1.4e+03| 1.1e+03| 1.6e+03|
Arp220          |CI2-1  | | 1.5e+03| 1.4e+03| 1.6e+03|
Arp220          |CO4-3  | | 3.2e+03| 2.8e+03| 3.5e+03|
Arp220          |CO5-4  | | 3.1e+03| 2.9e+03| 3.3e+03|
Arp220          |CO6-5  | | 3.4e+03| 3.2e+03| 3.6e+03|
Arp220          |CO7-6  | | 2.9e+03| 2.8e+03| 3.0e+03|
Arp220          |CO8-7  |X| 3.6e+03| 3.0e+03| 4.1e+03|
Arp220          |CO9-8  | | 2.3e+03| 2.0e+03| 2.6e+03|
Arp220          |CO10-9 | | 2.1e+03| 1.8e+03| 2.4e+03|
Arp220          |CO11-10| | 1.0e+03| 9.0e+02| 1.2e+03|
Arp220          |CO12-11| | 6.5e+02| 5.3e+02| 7.7e+02| 1.3e+03
Arp220          |CO13-12| | 3.6e+02| 1.9e+02| 5.3e+02| 1.1e+03
Arp220          |NII    |X| 2.2e+03| 1.7e+03| 2.7e+03|
NGC5990         |CI1-0  | | 4.1e+02| 1.8e+02| 6.8e+02| 1.0e+03
NGC5990         |CI2-1  | | 4.5e+02| 3.4e+02| 5.5e+02|
NGC5990         |CO4-3  | | 3.2e+02| 8.7e+01| 5.5e+02| 9.0e+02
NGC5990         |CO5-4  | | 7.3e+02| 5.5e+02| 9.2e+02|
NGC5990         |CO6-5  | | 4.8e+02| 3.6e+02| 5.9e+02|
NGC5990         |CO7-6  | | 3.2e+02| 2.2e+02| 4.2e+02|
NGC5990         |CO8-7  | | 3.8e+02| 2.3e+02| 5.4e+02|
NGC5990         |CO9-8  | | 1.5e+02| 3.1e+01| 3.1e+02| 5.6e+02
NGC5990         |CO10-9 | | 2.3e+02| 9.7e+01| 3.6e+02| 5.7e+02
NGC5990         |CO11-10| | 1.3e+02| 2.8e+01| 2.2e+02| 3.2e+02
NGC5990         |CO12-11| | 1.5e+02| 6.6e+01| 2.6e+02| 4.4e+02
NGC5990         |CO13-12| | 1.0e+02| 2.0e+01| 2.1e+02| 3.9e+02
NGC5990         |NII    | | 2.8e+03| 2.7e+03| 2.9e+03|
IRAS 15462-0450 |CI2-1  | | 3.5e+01| 7.5e+00| 6.8e+01| 1.1e+02
IRAS 15462-0450 |CO5-4  | | 1.1e+02| 2.6e+01| 2.5e+02| 4.2e+02
IRAS 15462-0450 |CO6-5  | | 7.9e+01| 2.9e+01| 1.3e+02| 2.2e+02
IRAS 15462-0450 |CO7-6  | | 1.4e+02| 1.0e+02| 1.8e+02|
IRAS 15462-0450 |CO8-7  | | 7.6e+01| 4.1e+01| 1.1e+02|
IRAS 15462-0450 |CO10-9 | | 7.2e+01| 3.2e+01| 1.1e+02| 1.7e+02
IRAS 15462-0450 |CO11-10| | 2.8e+01| 4.6e+00| 6.5e+01| 1.2e+02
IRAS 15462-0450 |CO12-11| | 3.9e+01| 1.0e+01| 7.9e+01| 1.2e+02
IRAS 15462-0450 |CO13-12| | 5.7e+01| 2.6e+01| 9.1e+01| 1.4e+02
IRAS 15462-0450 |NII    | | 1.1e+02| 7.6e+01| 1.5e+02|
3C 326          |CO5-4  | | 1.2e+02| 3.2e+01| 2.0e+02| 3.7e+02
3C 326          |CO7-6  | | 2.9e+01| 8.3e+00| 5.7e+01| 8.8e+01
3C 326          |CO8-7  | | 3.2e+01| 7.7e+00| 6.3e+01| 1.2e+02
3C 326          |CO9-8  | | 9.7e+01| 4.2e+01| 1.6e+02| 2.5e+02
3C 326          |CO10-9 | | 2.1e+01| 5.1e+00| 5.8e+01| 9.5e+01
3C 326          |CO11-10| | 4.2e+01| 1.3e+01| 7.1e+01| 1.2e+02
3C 326          |NII    | | 2.8e+01| 5.6e+00| 5.2e+01| 9.0e+01
PKS 1549-79     |CI2-1  | | 2.8e+01| 6.5e+00| 6.4e+01| 1.2e+02
PKS 1549-79     |CO5-4  | | 2.6e+02| 1.4e+02| 4.0e+02| 6.4e+02
PKS 1549-79     |CO6-5  | | 7.3e+01| 1.9e+01| 1.4e+02| 2.6e+02
PKS 1549-79     |CO7-6  | | 3.4e+01| 7.3e+00| 7.1e+01| 1.3e+02
PKS 1549-79     |CO10-9 | | 2.9e+01| 4.8e+00| 7.8e+01| 1.4e+02
PKS 1549-79     |CO11-10| | 3.1e+01| 7.8e+00| 6.4e+01| 1.0e+02
PKS 1549-79     |CO12-11| | 4.4e+01| 1.3e+01| 7.7e+01| 1.4e+02
PKS 1549-79     |CO13-12| | 3.6e+01| 9.5e+00| 7.0e+01| 1.3e+02
NGC6052         |CI1-0  | | 9.4e+02| 6.3e+02| 1.3e+03|
NGC6052         |CI2-1  | | 1.6e+02| 8.8e+01| 2.2e+02|
NGC6052         |CO4-3  | | 1.4e+03| 1.0e+03| 1.9e+03|
NGC6052         |CO5-4  | | 6.9e+02| 4.5e+02| 9.0e+02|
NGC6052         |CO6-5  | | 5.2e+02| 4.1e+02| 6.2e+02|
NGC6052         |CO7-6  | | 8.6e+01| 2.7e+01| 1.6e+02| 2.4e+02
NGC6052         |CO8-7  | | 1.2e+02| 5.3e+01| 1.8e+02| 2.6e+02
NGC6052         |CO9-8  | | 1.6e+02| 4.9e+01| 2.8e+02| 4.4e+02
NGC6052         |CO11-10| | 2.1e+02| 8.1e+01| 3.3e+02| 5.0e+02
NGC6052         |CO12-11| | 7.3e+01| 1.4e+01| 1.4e+02| 2.7e+02
NGC6052         |CO13-12| | 1.1e+02| 3.0e+01| 2.0e+02| 3.5e+02
NGC6052         |NII    | | 6.6e+02| 5.8e+02| 7.7e+02|
IRAS 16090-0139 |CI2-1  | | 1.5e+02| 1.1e+02| 2.0e+02|
IRAS 16090-0139 |CO5-4  | | 2.5e+02| 8.1e+01| 4.1e+02| 6.9e+02
IRAS 16090-0139 |CO6-5  | | 1.4e+02| 4.4e+01| 2.4e+02| 3.8e+02
IRAS 16090-0139 |CO7-6  | | 3.9e+02| 3.4e+02| 4.4e+02|
IRAS 16090-0139 |CO8-7  | | 3.6e+02| 3.2e+02| 4.0e+02|
IRAS 16090-0139 |CO10-9 | | 2.7e+02| 1.9e+02| 3.3e+02|
IRAS 16090-0139 |CO11-10| | 1.6e+02| 1.1e+02| 2.0e+02|
IRAS 16090-0139 |CO12-11| | 8.2e+01| 3.7e+01| 1.2e+02| 1.9e+02
IRAS 16090-0139 |CO13-12| | 9.7e+01| 6.1e+01| 1.3e+02|
IRAS 16090-0139 |NII    | | 4.9e+01| 1.6e+01| 7.8e+01| 1.4e+02
PG 1613+658     |CI2-1  | | 4.5e+01| 1.4e+01| 9.1e+01| 1.6e+02
PG 1613+658     |CO5-4  | | 8.2e+01| 1.1e+01| 2.1e+02| 4.5e+02
PG 1613+658     |CO6-5  | | 1.2e+02| 4.1e+01| 2.1e+02| 3.9e+02
PG 1613+658     |CO8-7  | | 2.6e+01| 5.2e+00| 5.1e+01| 1.1e+02
PG 1613+658     |CO10-9 | | 5.8e+01| 1.9e+01| 1.1e+02| 1.6e+02
PG 1613+658     |CO12-11| | 5.7e+01| 1.9e+01| 1.0e+02| 1.7e+02
PG 1613+658     |CO13-12| | 3.9e+01| 1.3e+01| 7.3e+01| 1.3e+02
PG 1613+658     |NII    | | 2.8e+01| 4.3e+00| 5.3e+01| 9.2e+01
CGCG052-037     |CI1-0  | | 7.3e+02| 4.8e+02| 9.5e+02|
CGCG052-037     |CI2-1  | | 4.1e+02| 3.6e+02| 4.6e+02|
CGCG052-037     |CO5-4  | | 7.6e+02| 5.8e+02| 9.5e+02|
CGCG052-037     |CO6-5  | | 5.7e+02| 4.9e+02| 6.4e+02|
CGCG052-037     |CO7-6  | | 3.4e+02| 2.8e+02| 3.8e+02|
CGCG052-037     |CO8-7  | | 2.4e+02| 2.0e+02| 3.0e+02|
CGCG052-037     |CO9-8  | | 6.6e+01| 2.0e+01| 1.3e+02| 2.2e+02
CGCG052-037     |CO10-9 | | 1.0e+02| 4.7e+01| 1.4e+02| 2.0e+02
CGCG052-037     |CO12-11| | 1.1e+02| 7.3e+01| 1.5e+02|
CGCG052-037     |NII    | | 1.2e+03| 1.2e+03| 1.3e+03|
NGC6156         |CI1-0  | | 4.4e+02| 2.0e+02| 7.2e+02| 1.1e+03
NGC6156         |CI2-1  | | 5.2e+02| 4.3e+02| 6.1e+02|
NGC6156         |CO4-3  | | 1.2e+03| 9.0e+02| 1.5e+03|
NGC6156         |CO5-4  | | 7.5e+02| 5.3e+02| 9.4e+02|
NGC6156         |CO6-5  | | 6.0e+02| 4.8e+02| 7.2e+02|
NGC6156         |CO7-6  | | 4.1e+02| 3.3e+02| 4.9e+02|
NGC6156         |CO8-7  | | 5.5e+02| 4.0e+02| 6.7e+02|
NGC6156         |CO9-8  | | 6.5e+02| 3.8e+02| 9.1e+02|
NGC6156         |CO10-9 | | 8.9e+01| 8.2e+00| 2.4e+02| 5.1e+02
NGC6156         |CO11-10| | 3.2e+02| 1.4e+02| 5.5e+02| 7.9e+02
NGC6156         |CO12-11| | 1.9e+02| 5.4e+01| 3.4e+02| 6.1e+02
NGC6156         |NII    | | 3.5e+03| 3.3e+03| 3.7e+03|
ESO069-IG006    |CI1-0  | | 8.2e+02| 5.7e+02| 1.1e+03|
ESO069-IG006    |CI2-1  | | 4.3e+02| 4.0e+02| 4.6e+02|
ESO069-IG006    |CO5-4  | | 1.1e+03| 9.3e+02| 1.2e+03|
ESO069-IG006    |CO6-5  | | 5.5e+02| 4.9e+02| 6.3e+02|
ESO069-IG006    |CO7-6  | | 2.9e+02| 2.5e+02| 3.2e+02|
ESO069-IG006    |CO8-7  | | 1.6e+02| 1.2e+02| 2.0e+02|
ESO069-IG006    |CO9-8  | | 6.9e+01| 2.2e+01| 1.3e+02| 2.3e+02
ESO069-IG006    |CO10-9 | | 8.7e+01| 3.6e+01| 1.3e+02| 1.8e+02
ESO069-IG006    |CO11-10| | 4.4e+01| 1.4e+01| 8.7e+01| 1.5e+02
ESO069-IG006    |CO12-11| | 3.9e+01| 1.1e+01| 7.6e+01| 1.2e+02
ESO069-IG006    |NII    |X| 2.0e+03| 1.9e+03| 2.0e+03|
IRASF16399-0937 |CI1-0  | | 1.2e+02| 3.6e+01| 2.2e+02| 4.5e+02
IRASF16399-0937 |CI2-1  | | 2.2e+02| 1.9e+02| 2.6e+02|
IRASF16399-0937 |CO5-4  | | 3.0e+02| 1.9e+02| 3.9e+02|
IRASF16399-0937 |CO6-5  | | 3.3e+02| 2.9e+02| 3.7e+02|
IRASF16399-0937 |CO7-6  | | 2.1e+02| 1.7e+02| 2.4e+02|
IRASF16399-0937 |CO8-7  | | 1.6e+02| 1.2e+02| 2.0e+02|
IRASF16399-0937 |CO9-8  | | 1.7e+02| 1.0e+02| 2.4e+02|
IRASF16399-0937 |CO10-9 | | 1.8e+02| 1.3e+02| 2.4e+02|
IRASF16399-0937 |CO11-10| | 7.1e+01| 2.0e+01| 1.2e+02| 2.2e+02
IRASF16399-0937 |CO12-11| | 9.4e+01| 4.3e+01| 1.4e+02| 2.2e+02
IRASF16399-0937 |CO13-12| | 7.4e+01| 3.1e+01| 1.1e+02| 1.8e+02
IRASF16399-0937 |NII    | | 8.9e+02| 8.4e+02| 9.3e+02|
NGC6240         |CI1-0  | | 2.0e+03| 1.7e+03| 2.2e+03|
NGC6240         |CI2-1  |X| 3.5e+03| 3.4e+03| 3.6e+03|
NGC6240         |CO4-3  | | 5.3e+03| 5.0e+03| 5.6e+03|
NGC6240         |CO5-4  | | 5.6e+03| 5.4e+03| 5.7e+03|
NGC6240         |CO6-5  |X| 6.8e+03| 6.7e+03| 7.0e+03|
NGC6240         |CO7-6  |X| 6.1e+03| 6.0e+03| 6.3e+03|
NGC6240         |CO8-7  |X| 5.1e+03| 5.0e+03| 5.3e+03|
NGC6240         |CO9-8  |X| 5.0e+03| 4.9e+03| 5.1e+03|
NGC6240         |CO10-9 |X| 4.5e+03| 4.4e+03| 4.6e+03|
NGC6240         |CO11-10|X| 3.4e+03| 3.3e+03| 3.4e+03|
NGC6240         |CO12-11|X| 2.6e+03| 2.6e+03| 2.7e+03|
NGC6240         |CO13-12|X| 2.2e+03| 2.2e+03| 2.3e+03|
NGC6240         |NII    |X| 3.8e+03| 3.7e+03| 3.9e+03|
IRASF16516-0948 |CI1-0  | | 1.4e+02| 5.2e+01| 2.1e+02| 4.1e+02
IRASF16516-0948 |CI2-1  | | 2.0e+02| 1.8e+02| 2.3e+02|
IRASF16516-0948 |CO5-4  | | 3.3e+02| 2.5e+02| 4.0e+02|
IRASF16516-0948 |CO6-5  | | 2.5e+02| 2.1e+02| 2.9e+02|
IRASF16516-0948 |CO7-6  | | 1.4e+02| 1.1e+02| 1.6e+02|
IRASF16516-0948 |CO8-7  | | 5.6e+01| 1.6e+01| 9.7e+01| 1.4e+02
IRASF16516-0948 |CO9-8  | | 1.8e+02| 1.0e+02| 2.5e+02|
IRASF16516-0948 |CO10-9 | | 7.4e+01| 2.9e+01| 1.3e+02| 2.0e+02
IRASF16516-0948 |CO12-11| | 6.3e+01| 1.9e+01| 1.2e+02| 1.9e+02
IRASF16516-0948 |CO13-12| | 7.6e+01| 2.8e+01| 1.3e+02| 2.0e+02
IRASF16516-0948 |NII    | | 9.0e+02| 8.5e+02| 9.6e+02|
NGC6286b        |CI1-0  | | 1.1e+02| 2.6e+01| 2.6e+02| 4.5e+02
NGC6286b        |CI2-1  | | 1.3e+02| 5.0e+01| 2.2e+02| 3.2e+02
NGC6286b        |CO5-4  | | 1.8e+02| 5.0e+01| 3.2e+02| 5.4e+02
NGC6286b        |CO6-5  | | 7.3e+01| 1.8e+01| 1.7e+02| 2.6e+02
NGC6286b        |CO7-6  | | 8.1e+01| 2.2e+01| 1.6e+02| 2.8e+02
NGC6286b        |CO8-7  | | 2.8e+02| 1.6e+02| 4.1e+02|
NGC6286b        |CO9-8  | | 1.4e+02| 3.6e+01| 2.7e+02| 4.8e+02
NGC6286b        |CO10-9 | | 1.7e+02| 6.8e+01| 2.6e+02| 4.6e+02
NGC6286b        |CO13-12| | 9.5e+01| 2.4e+01| 1.7e+02| 3.8e+02
NGC6286b        |NII    | | 6.1e+02| 4.9e+02| 7.2e+02|
NGC6286a        |CI1-0  | | 1.0e+03| 6.7e+02| 1.3e+03|
NGC6286a        |CI2-1  | | 7.4e+02| 6.5e+02| 8.3e+02|
NGC6286a        |CO5-4  | | 7.6e+02| 4.9e+02| 1.0e+03|
NGC6286a        |CO6-5  | | 5.0e+02| 3.7e+02| 6.0e+02|
NGC6286a        |CO7-6  | | 2.2e+02| 1.3e+02| 3.1e+02|
NGC6286a        |CO8-7  | | 3.0e+02| 1.8e+02| 4.3e+02|
NGC6286a        |CO9-8  | | 1.4e+02| 4.2e+01| 2.6e+02| 5.1e+02
NGC6286a        |CO11-10| | 1.2e+02| 3.7e+01| 2.2e+02| 4.0e+02
NGC6286a        |CO13-12| | 1.4e+02| 4.6e+01| 2.5e+02| 4.0e+02
NGC6286a        |NII    |X| 6.0e+03| 5.8e+03| 6.1e+03|
IRASF17138-1017 |CI2-1  | | 5.1e+02| 4.2e+02| 5.7e+02|
IRASF17138-1017 |CO4-3  | | 1.2e+03| 8.1e+02| 1.4e+03|
IRASF17138-1017 |CO5-4  | | 7.0e+02| 5.0e+02| 8.6e+02|
IRASF17138-1017 |CO6-5  | | 6.0e+02| 4.9e+02| 7.0e+02|
IRASF17138-1017 |CO7-6  | | 6.2e+02| 5.4e+02| 6.9e+02|
IRASF17138-1017 |CO8-7  | | 2.8e+02| 1.7e+02| 3.9e+02|
IRASF17138-1017 |CO9-8  | | 3.1e+02| 1.4e+02| 4.7e+02| 6.9e+02
IRASF17138-1017 |CO10-9 | | 3.0e+02| 2.0e+02| 3.9e+02|
IRASF17138-1017 |CO11-10| | 1.2e+02| 3.4e+01| 2.3e+02| 3.7e+02
IRASF17138-1017 |CO12-11| | 1.3e+02| 3.9e+01| 2.1e+02| 3.4e+02
IRASF17138-1017 |NII    | | 1.8e+03| 1.7e+03| 1.9e+03|
IRAS F17207-0014|CI1-0  | | 5.9e+02| 2.9e+02| 8.6e+02| 1.3e+03
IRAS F17207-0014|CI2-1  | | 7.3e+02| 6.5e+02| 7.9e+02|
IRAS F17207-0014|CO5-4  | | 1.2e+03| 1.0e+03| 1.3e+03|
IRAS F17207-0014|CO6-5  | | 1.3e+03| 1.2e+03| 1.4e+03|
IRAS F17207-0014|CO7-6  | | 1.2e+03| 1.1e+03| 1.3e+03|
IRAS F17207-0014|CO8-7  | | 1.1e+03| 9.8e+02| 1.1e+03|
IRAS F17207-0014|CO9-8  |X| 1.1e+03| 8.8e+02| 1.2e+03|
IRAS F17207-0014|CO10-9 |X| 1.4e+03| 1.3e+03| 1.6e+03|
IRAS F17207-0014|CO11-10|X| 7.4e+02| 6.1e+02| 8.7e+02|
IRAS F17207-0014|CO12-11|X| 5.1e+02| 3.9e+02| 6.4e+02|
IRAS F17207-0014|CO13-12|X| 3.1e+02| 2.1e+02| 4.1e+02|
IRAS F17207-0014|NII    |X| 1.1e+03| 9.8e+02| 1.2e+03|
ESO138-G027     |CI1-0  | | 1.6e+02| 3.7e+01| 4.2e+02| 7.9e+02
ESO138-G027     |CI2-1  | | 1.4e+02| 1.0e+02| 2.0e+02|
ESO138-G027     |CO5-4  | | 5.0e+02| 3.2e+02| 6.4e+02|
ESO138-G027     |CO6-5  | | 1.8e+02| 1.0e+02| 2.5e+02|
ESO138-G027     |CO7-6  | | 2.3e+02| 1.9e+02| 2.8e+02|
ESO138-G027     |CO8-7  | | 1.5e+02| 8.2e+01| 2.1e+02|
ESO138-G027     |CO9-8  | | 1.1e+02| 2.6e+01| 2.0e+02| 3.9e+02
ESO138-G027     |CO10-9 | | 1.2e+02| 5.7e+01| 2.0e+02| 3.2e+02
ESO138-G027     |CO11-10| | 1.6e+02| 8.2e+01| 2.4e+02| 4.0e+02
ESO138-G027     |CO12-11| | 1.4e+02| 7.3e+01| 2.2e+02| 3.0e+02
ESO138-G027     |CO13-12| | 1.5e+02| 7.3e+01| 2.2e+02| 3.2e+02
ESO138-G027     |NII    | | 1.2e+03| 1.2e+03| 1.3e+03|
UGC11041        |CI1-0  | | 2.9e+02| 5.9e+01| 6.4e+02| 1.0e+03
UGC11041        |CI2-1  | | 4.0e+02| 3.5e+02| 4.7e+02|
UGC11041        |CO4-3  | | 4.4e+02| 1.7e+02| 7.8e+02| 1.7e+03
UGC11041        |CO5-4  | | 3.6e+02| 1.5e+02| 5.6e+02| 8.6e+02
UGC11041        |CO6-5  | | 2.6e+02| 1.8e+02| 3.5e+02|
UGC11041        |CO7-6  | | 2.1e+02| 1.5e+02| 2.7e+02|
UGC11041        |CO9-8  | | 2.4e+02| 1.5e+02| 3.3e+02| 4.6e+02
UGC11041        |CO13-12| | 6.7e+01| 1.6e+01| 1.4e+02| 2.4e+02
UGC11041        |NII    | | 2.0e+03| 1.9e+03| 2.1e+03|
IRAS17578-0400  |CI1-0  | | 2.3e+02| 4.7e+01| 5.0e+02| 8.2e+02
IRAS17578-0400  |CI2-1  | | 3.9e+02| 3.2e+02| 4.7e+02|
IRAS17578-0400  |CO4-3  | | 4.4e+02| 2.0e+02| 7.6e+02| 1.1e+03
IRAS17578-0400  |CO5-4  | | 4.8e+02| 3.0e+02| 6.8e+02|
IRAS17578-0400  |CO6-5  | | 7.4e+02| 6.4e+02| 8.1e+02|
IRAS17578-0400  |CO7-6  | | 5.6e+02| 4.8e+02| 6.3e+02|
IRAS17578-0400  |CO8-7  | | 5.1e+02| 3.9e+02| 6.0e+02|
IRAS17578-0400  |CO9-8  | | 7.4e+02| 6.2e+02| 8.5e+02|
IRAS17578-0400  |CO10-9 | | 4.2e+02| 3.1e+02| 5.3e+02|
IRAS17578-0400  |CO11-10| | 2.7e+02| 1.5e+02| 3.8e+02| 5.6e+02
IRAS17578-0400  |CO12-11| | 1.4e+02| 5.4e+01| 2.2e+02| 3.6e+02
IRAS17578-0400  |NII    | | 9.6e+02| 8.6e+02| 1.1e+03|
NGC6621         |CI1-0  | | 6.5e+02| 3.0e+02| 9.3e+02| 1.5e+03
NGC6621         |CI2-1  | | 5.0e+02| 4.2e+02| 5.7e+02|
NGC6621         |CO5-4  | | 9.1e+02| 6.5e+02| 1.2e+03|
NGC6621         |CO6-5  | | 9.1e+02| 8.0e+02| 1.0e+03|
NGC6621         |CO7-6  | | 2.9e+02| 2.2e+02| 3.6e+02|
NGC6621         |CO9-8  | | 1.0e+02| 2.6e+01| 1.8e+02| 4.2e+02
NGC6621         |CO10-9 | | 1.7e+02| 7.4e+01| 2.6e+02| 3.9e+02
NGC6621         |CO13-12| | 7.5e+01| 2.2e+01| 1.5e+02| 2.4e+02
NGC6621         |NII    | | 1.4e+03| 1.3e+03| 1.5e+03|
IC4687          |CI1-0  | | 3.2e+02| 2.2e+02| 4.1e+02|
IC4687          |CI2-1  | | 5.5e+02| 5.1e+02| 5.8e+02|
IC4687          |CO4-3  | | 6.1e+02| 5.0e+02| 7.2e+02|
IC4687          |CO5-4  | | 6.5e+02| 5.9e+02| 7.2e+02|
IC4687          |CO6-5  | | 7.3e+02| 6.8e+02| 7.7e+02|
IC4687          |CO7-6  | | 5.4e+02| 5.0e+02| 5.7e+02|
IC4687          |CO8-7  | | 3.7e+02| 3.2e+02| 4.1e+02|
IC4687          |CO9-8  | | 1.5e+02| 9.8e+01| 2.0e+02|
IC4687          |CO10-9 | | 1.5e+02| 1.2e+02| 1.9e+02|
IC4687          |CO11-10| | 2.1e+01| 3.0e+00| 5.1e+01| 1.2e+02
IC4687          |CO12-11| | 6.1e+01| 3.5e+01| 9.3e+01| 1.3e+02
IC4687          |CO13-12| | 3.3e+01| 6.0e+00| 7.2e+01| 1.4e+02
IC4687          |NII    | | 2.3e+03| 2.2e+03| 2.3e+03|
IRAS F18293-3413|CI1-0  | | 2.3e+03| 2.1e+03| 2.5e+03|
IRAS F18293-3413|CI2-1  | | 2.3e+03| 2.2e+03| 2.3e+03|
IRAS F18293-3413|CO4-3  | | 3.4e+03| 3.2e+03| 3.6e+03|
IRAS F18293-3413|CO5-4  | | 3.2e+03| 3.1e+03| 3.4e+03|
IRAS F18293-3413|CO6-5  | | 2.8e+03| 2.8e+03| 2.9e+03|
IRAS F18293-3413|CO7-6  | | 1.9e+03| 1.9e+03| 2.0e+03|
IRAS F18293-3413|CO8-7  | | 1.1e+03| 1.0e+03| 1.2e+03|
IRAS F18293-3413|CO9-8  | | 7.9e+02| 6.9e+02| 8.9e+02|
IRAS F18293-3413|CO10-9 | | 4.2e+02| 3.5e+02| 4.9e+02|
IRAS F18293-3413|CO11-10| | 2.2e+02| 1.4e+02| 2.9e+02|
IRAS F18293-3413|CO12-11| | 1.4e+02| 7.8e+01| 2.3e+02| 3.0e+02
IRAS F18293-3413|CO13-12| | 1.5e+02| 6.4e+01| 2.4e+02| 3.4e+02
IRAS F18293-3413|NII    |X| 5.7e+03| 5.6e+03| 5.8e+03|
IC4734          |CI1-0  | | 4.0e+02| 1.5e+02| 7.7e+02| 1.2e+03
IC4734          |CI2-1  | | 5.8e+02| 4.9e+02| 6.7e+02|
IC4734          |CO5-4  | | 1.4e+03| 1.1e+03| 1.6e+03|
IC4734          |CO6-5  | | 1.1e+03| 9.0e+02| 1.2e+03|
IC4734          |CO7-6  | | 6.6e+02| 5.6e+02| 7.6e+02|
IC4734          |CO8-7  | | 5.9e+02| 4.7e+02| 7.0e+02|
IC4734          |CO9-8  | | 4.8e+02| 3.4e+02| 6.1e+02|
IC4734          |CO10-9 | | 3.5e+02| 2.4e+02| 4.4e+02|
IC4734          |CO11-10| | 2.7e+02| 1.5e+02| 4.0e+02| 5.6e+02
IC4734          |CO12-11| | 1.5e+02| 6.3e+01| 2.4e+02| 3.4e+02
IC4734          |CO13-12| | 2.2e+02| 9.8e+01| 3.5e+02| 5.1e+02
IC4734          |NII    | | 1.2e+03| 1.1e+03| 1.3e+03|
NGC6701         |CI1-0  | | 1.2e+03| 8.0e+02| 1.6e+03|
NGC6701         |CI2-1  | | 7.6e+02| 6.7e+02| 8.4e+02|
NGC6701         |CO4-3  | | 1.0e+03| 6.4e+02| 1.4e+03| 2.0e+03
NGC6701         |CO5-4  | | 1.4e+03| 1.1e+03| 1.7e+03|
NGC6701         |CO6-5  | | 9.5e+02| 8.2e+02| 1.1e+03|
NGC6701         |CO7-6  | | 5.8e+02| 4.8e+02| 6.5e+02|
NGC6701         |CO8-7  | | 5.1e+02| 3.9e+02| 6.4e+02|
NGC6701         |CO9-8  | | 5.2e+02| 3.4e+02| 6.6e+02|
NGC6701         |CO10-9 | | 4.8e+02| 3.2e+02| 6.2e+02|
NGC6701         |CO11-10| | 1.5e+02| 3.0e+01| 2.7e+02| 4.6e+02
NGC6701         |CO12-11| | 1.8e+02| 6.6e+01| 2.9e+02| 4.5e+02
NGC6701         |CO13-12| | 2.4e+02| 1.1e+02| 3.9e+02| 5.6e+02
NGC6701         |NII    | | 1.9e+03| 1.7e+03| 2.0e+03|
IRAS 19254-7245 |CI2-1  | | 2.9e+02| 2.4e+02| 3.4e+02|
IRAS 19254-7245 |CO7-6  | | 3.7e+02| 3.2e+02| 4.2e+02|
IRAS 19254-7245 |CO8-7  | | 2.2e+02| 1.5e+02| 2.8e+02|
IRAS 19254-7245 |CO9-8  | | 3.0e+02| 2.2e+02| 3.7e+02|
IRAS 19254-7245 |CO10-9 | | 1.8e+02| 1.3e+02| 2.4e+02|
IRAS 19254-7245 |CO11-10| | 1.1e+02| 5.3e+01| 1.6e+02| 2.3e+02
IRAS 19254-7245 |CO12-11| | 5.1e+01| 1.9e+01| 9.2e+01| 1.5e+02
IRAS 19254-7245 |CO13-12| | 1.0e+02| 5.9e+01| 1.5e+02|
IRAS 19254-7245 |NII    |X| 4.2e+02| 3.5e+02| 5.0e+02|
IRAS 19297-0406 |CI1-0  | | 3.2e+02| 1.4e+02| 4.7e+02| 8.0e+02
IRAS 19297-0406 |CI2-1  | | 1.3e+02| 9.2e+01| 1.7e+02|
IRAS 19297-0406 |CO5-4  | | 1.9e+02| 7.8e+01| 3.6e+02| 5.8e+02
IRAS 19297-0406 |CO6-5  | | 1.5e+02| 7.7e+01| 2.2e+02| 3.3e+02
IRAS 19297-0406 |CO7-6  | | 1.6e+02| 1.2e+02| 1.9e+02|
IRAS 19297-0406 |CO8-7  | | 1.7e+02| 1.4e+02| 2.0e+02|
IRAS 19297-0406 |CO9-8  | | 1.1e+02| 3.1e+01| 1.8e+02| 2.5e+02
IRAS 19297-0406 |CO10-9 | | 1.8e+02| 1.1e+02| 2.4e+02|
IRAS 19297-0406 |CO11-10| | 1.0e+02| 4.3e+01| 1.7e+02| 2.6e+02
IRAS 19297-0406 |CO12-11| | 4.1e+01| 7.7e+00| 9.6e+01| 2.0e+02
IRAS 19297-0406 |CO13-12| | 7.6e+01| 2.1e+01| 1.3e+02| 2.1e+02
IRAS 19297-0406 |NII    | | 1.1e+02| 5.7e+01| 1.6e+02|
ESO339-G011     |CI1-0  | | 4.0e+02| 1.6e+02| 6.4e+02| 1.1e+03
ESO339-G011     |CI2-1  | | 3.2e+02| 2.6e+02| 3.8e+02|
ESO339-G011     |CO5-4  | | 3.7e+02| 2.0e+02| 5.5e+02| 8.1e+02
ESO339-G011     |CO6-5  | | 2.0e+02| 1.1e+02| 2.8e+02| 4.2e+02
ESO339-G011     |CO7-6  | | 1.9e+02| 1.3e+02| 2.4e+02|
ESO339-G011     |CO8-7  | | 1.4e+02| 5.3e+01| 2.3e+02| 3.9e+02
ESO339-G011     |CO9-8  | | 1.6e+02| 6.1e+01| 2.7e+02| 5.4e+02
ESO339-G011     |CO10-9 | | 1.5e+02| 6.0e+01| 2.5e+02| 4.0e+02
ESO339-G011     |CO11-10| | 1.8e+02| 7.3e+01| 3.0e+02| 4.1e+02
ESO339-G011     |CO12-11| | 9.8e+01| 2.4e+01| 1.6e+02| 2.9e+02
ESO339-G011     |NII    | | 1.3e+03| 1.2e+03| 1.4e+03|
3C 405          |CI1-0  | | 1.8e+02| 7.0e+01| 2.7e+02| 5.6e+02
3C 405          |CI2-1  | | 2.4e+02| 2.0e+02| 2.7e+02|
3C 405          |CO5-4  | | 1.4e+02| 5.2e+01| 2.8e+02| 4.3e+02
3C 405          |CO6-5  | | 9.3e+01| 3.4e+01| 1.4e+02| 2.2e+02
3C 405          |CO7-6  | | 3.7e+01| 9.6e+00| 6.7e+01| 1.3e+02
3C 405          |CO9-8  | | 1.0e+02| 4.6e+01| 1.7e+02| 2.4e+02
3C 405          |CO11-10| | 4.4e+01| 1.6e+01| 8.7e+01| 1.4e+02
3C 405          |CO13-12| | 5.2e+01| 2.1e+01| 9.2e+01| 1.4e+02
3C 405          |NII    | | 3.4e+02| 3.1e+02| 3.8e+02|
IRAS 20087-0308 |CI2-1  | | 2.0e+02| 1.5e+02| 2.4e+02|
IRAS 20087-0308 |CO5-4  | | 4.8e+02| 2.6e+02| 6.3e+02|
IRAS 20087-0308 |CO6-5  | | 1.4e+02| 7.0e+01| 2.2e+02| 3.2e+02
IRAS 20087-0308 |CO7-6  | | 3.1e+02| 2.7e+02| 3.5e+02|
IRAS 20087-0308 |CO8-7  | | 1.9e+02| 1.5e+02| 2.3e+02|
IRAS 20087-0308 |CO10-9 | | 2.0e+02| 1.4e+02| 2.5e+02|
IRAS 20087-0308 |CO11-10| | 8.3e+01| 3.6e+01| 1.3e+02| 1.9e+02
IRAS 20087-0308 |CO12-11| | 6.8e+01| 2.2e+01| 1.2e+02| 1.9e+02
IRAS 20087-0308 |CO13-12| | 9.6e+01| 5.7e+01| 1.3e+02|
IRAS 20087-0308 |NII    | | 1.3e+02| 8.3e+01| 1.7e+02|
IRAS 20100-4156 |CI2-1  | | 1.6e+02| 1.1e+02| 2.0e+02|
IRAS 20100-4156 |CO5-4  | | 3.3e+02| 1.7e+02| 4.7e+02|
IRAS 20100-4156 |CO6-5  | | 8.2e+01| 1.7e+01| 1.7e+02| 3.2e+02
IRAS 20100-4156 |CO7-6  | | 1.7e+02| 1.2e+02| 2.1e+02|
IRAS 20100-4156 |CO8-7  | | 2.0e+02| 1.5e+02| 2.4e+02|
IRAS 20100-4156 |CO10-9 | | 2.2e+02| 1.6e+02| 2.7e+02|
IRAS 20100-4156 |CO11-10| | 7.2e+01| 3.1e+01| 1.2e+02| 1.7e+02
IRAS 20100-4156 |CO12-11| | 9.1e+01| 3.7e+01| 1.4e+02| 2.0e+02
IRAS 20100-4156 |CO13-12| | 5.6e+01| 2.3e+01| 9.1e+01| 1.4e+02
IRAS 20100-4156 |NII    | | 1.7e+02| 1.3e+02| 2.1e+02|
MCG+04-48-002a  |CI1-0  | | 5.1e+02| 1.5e+02| 9.2e+02| 1.6e+03
MCG+04-48-002a  |CI2-1  | | 5.0e+02| 4.1e+02| 5.9e+02|
MCG+04-48-002a  |CO5-4  | | 8.1e+02| 5.4e+02| 1.0e+03|
MCG+04-48-002a  |CO6-5  | | 3.2e+02| 1.9e+02| 4.8e+02| 6.2e+02
MCG+04-48-002a  |CO7-6  | | 3.5e+02| 2.8e+02| 4.4e+02|
MCG+04-48-002a  |CO8-7  | | 3.3e+02| 2.0e+02| 4.6e+02| 6.6e+02
MCG+04-48-002a  |CO10-9 | | 1.2e+02| 3.2e+01| 2.3e+02| 4.2e+02
MCG+04-48-002a  |CO11-10| | 2.0e+02| 8.0e+01| 3.2e+02| 4.7e+02
MCG+04-48-002a  |CO12-11| | 3.6e+01| 4.8e+00| 1.1e+02| 2.4e+02
MCG+04-48-002a  |NII    |X| 3.1e+03| 2.9e+03| 3.2e+03|
NGC6926         |CI1-0  | | 4.6e+02| 2.2e+02| 7.0e+02| 1.1e+03
NGC6926         |CI2-1  | | 3.3e+02| 2.7e+02| 4.0e+02|
NGC6926         |CO5-4  | | 4.9e+02| 3.4e+02| 6.5e+02|
NGC6926         |CO6-5  | | 7.3e+01| 1.8e+01| 1.5e+02| 2.5e+02
NGC6926         |CO7-6  | | 1.3e+02| 8.7e+01| 2.0e+02|
NGC6926         |CO9-8  | | 1.1e+02| 2.0e+01| 2.5e+02| 4.2e+02
NGC6926         |CO10-9 | | 2.0e+02| 6.6e+01| 3.4e+02| 6.1e+02
NGC6926         |CO11-10| | 2.0e+02| 6.8e+01| 3.4e+02| 5.7e+02
NGC6926         |CO12-11| | 1.5e+02| 4.4e+01| 3.1e+02| 4.9e+02
NGC6926         |CO13-12| | 2.5e+02| 1.0e+02| 3.9e+02| 6.5e+02
NGC6926         |NII    | | 1.3e+03| 1.1e+03| 1.4e+03|
NGC6946         |CI1-0  | | 3.8e+03| 3.4e+03| 4.0e+03|
NGC6946         |CI2-1  | | 3.0e+03| 2.9e+03| 3.2e+03|
NGC6946         |CO4-3  | | 8.7e+03| 8.3e+03| 9.0e+03|
NGC6946         |CO5-4  | | 7.0e+03| 6.8e+03| 7.2e+03|
NGC6946         |CO6-5  | | 4.8e+03| 4.7e+03| 5.0e+03|
NGC6946         |CO7-6  | | 3.3e+03| 3.2e+03| 3.4e+03|
NGC6946         |CO8-7  | | 2.1e+03| 1.9e+03| 2.3e+03|
NGC6946         |CO9-8  | | 2.3e+03| 2.0e+03| 2.5e+03|
NGC6946         |CO10-9 | | 1.4e+03| 1.1e+03| 1.6e+03|
NGC6946         |CO11-10| | 1.2e+03| 9.0e+02| 1.5e+03|
NGC6946         |CO12-11| | 3.4e+02| 9.4e+01| 5.7e+02| 9.1e+02
NGC6946         |NII    | | 9.7e+03| 9.3e+03| 1.0e+04|
NGC6946_05      |CI1-0  | | 1.4e+02| 3.4e+01| 2.3e+02| 4.0e+02
NGC6946_05      |CI2-1  | | 2.2e+02| 1.4e+02| 2.7e+02|
NGC6946_05      |CO4-3  | | 6.5e+02| 4.5e+02| 8.3e+02|
NGC6946_05      |CO5-4  | | 1.6e+02| 5.0e+01| 3.0e+02| 4.7e+02
NGC6946_05      |CO6-5  | | 1.7e+02| 9.6e+01| 2.4e+02| 3.6e+02
NGC6946_05      |CO7-6  | | 2.0e+02| 1.3e+02| 2.5e+02|
NGC6946_05      |CO8-7  | | 9.1e+01| 2.3e+01| 1.5e+02| 2.3e+02
NGC6946_05      |CO9-8  | | 2.9e+02| 1.5e+02| 4.5e+02| 6.5e+02
NGC6946_05      |CO10-9 | | 6.0e+01| 7.6e+00| 1.6e+02| 3.7e+02
NGC6946_05      |CO12-11| | 1.3e+02| 3.6e+01| 2.7e+02| 4.8e+02
NGC6946_05      |CO13-12| | 1.8e+02| 4.5e+01| 3.4e+02| 6.0e+02
NGC6946_05      |NII    | | 5.3e+03| 5.2e+03| 5.5e+03|
IRAS 20414-1651 |CI2-1  | | 1.2e+02| 8.0e+01| 1.5e+02|
IRAS 20414-1651 |CO5-4  | | 1.4e+02| 3.4e+01| 2.6e+02| 4.3e+02
IRAS 20414-1651 |CO6-5  | | 6.9e+01| 2.1e+01| 1.2e+02| 2.0e+02
IRAS 20414-1651 |CO7-6  | | 7.2e+01| 3.5e+01| 1.1e+02| 1.9e+02
IRAS 20414-1651 |CO8-7  | | 1.4e+02| 9.1e+01| 1.8e+02|
IRAS 20414-1651 |CO9-8  | | 1.0e+02| 3.6e+01| 1.8e+02| 2.6e+02
IRAS 20414-1651 |CO10-9 | | 9.9e+01| 4.8e+01| 1.5e+02| 2.1e+02
IRAS 20414-1651 |CO11-10| | 3.3e+01| 1.1e+01| 7.3e+01| 1.4e+02
IRAS 20414-1651 |CO12-11| | 1.0e+02| 6.4e+01| 1.4e+02|
IRAS 20414-1651 |CO13-12| | 4.5e+01| 1.8e+01| 7.7e+01| 1.2e+02
IRAS 20414-1651 |NII    | | 4.9e+01| 1.5e+01| 8.8e+01| 1.4e+02
3C 424          |CI2-1  | | 2.8e+01| 5.9e+00| 5.6e+01| 1.1e+02
3C 424          |CO5-4  | | 1.4e+02| 4.0e+01| 2.6e+02| 5.0e+02
3C 424          |CO6-5  | | 4.0e+01| 6.2e+00| 1.1e+02| 2.2e+02
3C 424          |CO8-7  | | 2.9e+01| 6.4e+00| 5.6e+01| 9.8e+01
3C 424          |CO10-9 | | 2.1e+01| 3.4e+00| 4.8e+01| 1.2e+02
3C 424          |CO11-10| | 5.7e+01| 2.8e+01| 1.0e+02| 1.5e+02
3C 424          |CO12-11| | 2.9e+01| 8.9e+00| 7.7e+01| 1.3e+02
3C 424          |CO13-12| | 1.9e+01| 2.5e+00| 3.8e+01| 8.9e+01
3C 424          |NII    | | 3.8e+01| 1.1e+01| 7.0e+01| 1.2e+02
IC 5063         |CI1-0  | | 4.7e+02| 1.3e+02| 8.9e+02| 1.4e+03
IC 5063         |CI2-1  | | 2.8e+02| 2.0e+02| 3.6e+02|
IC 5063         |CO5-4  | | 4.7e+02| 2.3e+02| 7.8e+02| 1.2e+03
IC 5063         |CO6-5  | | 2.1e+02| 8.5e+01| 3.3e+02| 5.0e+02
IC 5063         |CO7-6  | | 3.3e+02| 2.3e+02| 4.2e+02|
IC 5063         |CO8-7  | | 1.2e+02| 4.5e+01| 2.2e+02| 4.9e+02
IC 5063         |CO9-8  | | 1.6e+02| 4.1e+01| 3.0e+02| 5.6e+02
IC 5063         |CO10-9 | | 1.6e+02| 4.6e+01| 3.4e+02| 5.5e+02
IC 5063         |CO12-11| | 1.8e+02| 7.3e+01| 3.0e+02| 4.4e+02
IC 5063         |CO13-12| | 1.6e+02| 4.8e+01| 2.8e+02| 4.4e+02
IC 5063         |NII    | | 3.1e+02| 1.7e+02| 4.6e+02|
CGCG448-020     |CI1-0  | | 2.8e+02| 7.3e+01| 6.0e+02| 8.1e+02
CGCG448-020     |CI2-1  | | 3.1e+02| 2.3e+02| 3.9e+02|
CGCG448-020     |CO5-4  | | 4.9e+02| 2.2e+02| 7.4e+02|
CGCG448-020     |CO6-5  | | 3.2e+02| 1.8e+02| 4.3e+02|
CGCG448-020     |CO7-6  | | 3.7e+02| 3.0e+02| 4.6e+02|
CGCG448-020     |CO8-7  | | 3.8e+02| 2.8e+02| 4.8e+02|
CGCG448-020     |CO9-8  | | 4.0e+02| 2.5e+02| 5.5e+02|
CGCG448-020     |CO10-9 | | 4.5e+02| 3.6e+02| 5.5e+02|
CGCG448-020     |CO11-10| | 3.3e+02| 2.1e+02| 4.6e+02|
CGCG448-020     |CO12-11| | 5.7e+02| 4.6e+02| 6.7e+02|
CGCG448-020     |CO13-12| | 2.2e+02| 1.3e+02| 3.2e+02| 4.6e+02
CGCG448-020     |NII    | | 4.0e+02| 3.0e+02| 4.9e+02|
ESO286-IG019    |CI1-0  | | 1.9e+02| 5.0e+01| 3.9e+02| 7.5e+02
ESO286-IG019    |CI2-1  | | 2.4e+02| 1.8e+02| 2.9e+02|
ESO286-IG019    |CO5-4  | | 7.9e+02| 6.2e+02| 9.6e+02|
ESO286-IG019    |CO6-5  | | 5.4e+02| 4.6e+02| 6.2e+02|
ESO286-IG019    |CO7-6  | | 7.0e+02| 6.4e+02| 7.4e+02|
ESO286-IG019    |CO8-7  | | 7.0e+02| 6.4e+02| 7.6e+02|
ESO286-IG019    |CO9-8  | | 4.3e+02| 3.3e+02| 5.0e+02|
ESO286-IG019    |CO10-9 | | 5.7e+02| 5.1e+02| 6.2e+02|
ESO286-IG019    |CO11-10| | 4.7e+02| 4.1e+02| 5.3e+02|
ESO286-IG019    |CO12-11| | 3.6e+02| 3.1e+02| 4.0e+02|
ESO286-IG019    |CO13-12| | 2.8e+02| 2.3e+02| 3.3e+02|
ESO286-IG019    |NII    | | 1.5e+02| 9.3e+01| 2.0e+02|
ESO286-G035     |CI1-0  | | 1.0e+03| 6.4e+02| 1.3e+03|
ESO286-G035     |CI2-1  | | 2.9e+02| 2.2e+02| 3.5e+02|
ESO286-G035     |CO4-3  | | 1.7e+03| 1.4e+03| 2.1e+03|
ESO286-G035     |CO5-4  | | 8.2e+02| 6.0e+02| 1.0e+03|
ESO286-G035     |CO6-5  | | 6.3e+02| 5.3e+02| 7.2e+02|
ESO286-G035     |CO7-6  | | 2.7e+02| 2.0e+02| 3.3e+02|
ESO286-G035     |CO8-7  | | 1.4e+02| 6.7e+01| 2.4e+02| 3.8e+02
ESO286-G035     |CO9-8  | | 1.7e+02| 5.8e+01| 2.7e+02| 4.1e+02
ESO286-G035     |CO10-9 | | 8.6e+01| 2.4e+01| 1.5e+02| 2.4e+02
ESO286-G035     |CO11-10| | 1.1e+02| 4.1e+01| 1.8e+02| 3.2e+02
ESO286-G035     |CO13-12| | 5.8e+01| 1.5e+01| 1.4e+02| 2.2e+02
ESO286-G035     |NII    | | 1.7e+03| 1.6e+03| 1.8e+03|
3C 433          |CI2-1  | | 6.3e+01| 2.5e+01| 1.0e+02| 1.6e+02
3C 433          |CO5-4  | | 1.4e+02| 4.2e+01| 2.4e+02| 4.5e+02
3C 433          |CO6-5  | | 9.9e+01| 2.6e+01| 1.7e+02| 2.7e+02
3C 433          |CO7-6  | | 4.4e+01| 1.2e+01| 7.8e+01| 1.3e+02
3C 433          |CO8-7  | | 3.4e+01| 6.6e+00| 6.2e+01| 1.2e+02
3C 433          |CO10-9 | | 3.0e+01| 5.5e+00| 4.8e+01| 9.0e+01
3C 433          |CO11-10| | 4.2e+01| 1.2e+01| 7.8e+01| 1.2e+02
3C 433          |CO12-11| | 3.1e+01| 5.9e+00| 6.6e+01| 1.1e+02
3C 433          |NII    | | 2.7e+01| 7.2e+00| 5.9e+01| 1.1e+02
NGC7130         |CI1-0  | | 8.4e+02| 5.5e+02| 1.1e+03|
NGC7130         |CI2-1  | | 1.0e+03| 9.4e+02| 1.0e+03|
NGC7130         |CO4-3  | | 2.3e+03| 1.9e+03| 2.6e+03|
NGC7130         |CO5-4  | | 1.8e+03| 1.6e+03| 2.0e+03|
NGC7130         |CO6-5  | | 1.3e+03| 1.2e+03| 1.4e+03|
NGC7130         |CO7-6  | | 9.9e+02| 9.5e+02| 1.0e+03|
NGC7130         |CO8-7  | | 6.5e+02| 5.9e+02| 7.1e+02|
NGC7130         |CO9-8  | | 7.0e+02| 6.2e+02| 7.8e+02|
NGC7130         |CO10-9 | | 4.8e+02| 4.0e+02| 5.5e+02|
NGC7130         |CO11-10| | 3.4e+02| 2.6e+02| 4.0e+02|
NGC7130         |CO12-11| | 2.3e+02| 1.7e+02| 3.0e+02|
NGC7130         |CO13-12| | 1.4e+02| 6.2e+01| 2.3e+02| 3.3e+02
NGC7130         |NII    | | 2.9e+03| 2.8e+03| 2.9e+03|
NGC7172         |CI1-0  | | 1.0e+03| 6.6e+02| 1.4e+03|
NGC7172         |CI2-1  | | 7.8e+02| 7.1e+02| 8.6e+02|
NGC7172         |CO4-3  | | 6.4e+02| 2.4e+02| 1.1e+03| 2.0e+03
NGC7172         |CO5-4  | | 2.5e+02| 4.5e+01| 5.2e+02| 8.0e+02
NGC7172         |CO6-5  | | 4.7e+02| 3.6e+02| 5.7e+02|
NGC7172         |CO7-6  | | 7.2e+01| 1.9e+01| 1.4e+02| 2.4e+02
NGC7172         |CO8-7  | | 1.2e+02| 4.8e+01| 2.0e+02| 3.4e+02
NGC7172         |CO9-8  | | 8.8e+01| 2.7e+01| 1.6e+02| 2.8e+02
NGC7172         |CO11-10| | 8.2e+01| 3.0e+01| 1.6e+02| 2.8e+02
NGC7172         |CO13-12| | 1.1e+02| 4.2e+01| 1.9e+02| 2.9e+02
NGC7172         |NII    |X| 4.5e+03| 4.4e+03| 4.6e+03|
ESO467-G027     |CI1-0  | | 5.9e+02| 2.1e+02| 1.0e+03| 1.5e+03
ESO467-G027     |CI2-1  | | 3.5e+02| 2.9e+02| 4.1e+02|
ESO467-G027     |CO5-4  | | 4.0e+02| 1.5e+02| 7.0e+02| 1.2e+03
ESO467-G027     |CO6-5  | | 1.1e+02| 2.6e+01| 2.3e+02| 3.4e+02
ESO467-G027     |CO7-6  | | 5.4e+01| 7.4e+00| 1.1e+02| 1.9e+02
ESO467-G027     |CO8-7  | | 6.9e+01| 2.1e+01| 1.2e+02| 2.5e+02
ESO467-G027     |CO9-8  | | 1.3e+02| 4.0e+01| 2.2e+02| 3.8e+02
ESO467-G027     |CO10-9 | | 1.7e+02| 6.9e+01| 2.8e+02| 4.6e+02
ESO467-G027     |CO12-11| | 1.3e+02| 3.9e+01| 2.2e+02| 3.1e+02
ESO467-G027     |NII    | | 2.9e+03| 2.8e+03| 3.0e+03|
IC5179          |CI1-0  | | 8.5e+02| 6.2e+02| 1.1e+03|
IC5179          |CI2-1  | | 7.6e+02| 6.5e+02| 8.6e+02|
IC5179          |CO4-3  | | 6.6e+02| 3.4e+02| 1.0e+03| 1.4e+03
IC5179          |CO5-4  | | 7.2e+02| 4.8e+02| 9.3e+02|
IC5179          |CO6-5  | | 6.7e+02| 5.4e+02| 7.9e+02|
IC5179          |CO7-6  | | 4.1e+02| 3.0e+02| 5.2e+02|
IC5179          |CO8-7  | | 2.4e+02| 1.0e+02| 3.9e+02| 6.4e+02
IC5179          |CO9-8  | | 2.0e+02| 5.6e+01| 3.6e+02| 5.9e+02
IC5179          |CO12-11| | 1.3e+02| 2.5e+01| 2.7e+02| 4.7e+02
IC5179          |NII    | | 6.5e+03| 6.4e+03| 6.7e+03|
NGC7331         |CI1-0  | | 9.1e+02| 6.2e+02| 1.2e+03|
NGC7331         |CI2-1  | | 7.1e+02| 6.4e+02| 7.8e+02|
NGC7331         |CO4-3  | | 1.6e+03| 1.3e+03| 1.8e+03|
NGC7331         |CO5-4  | | 6.6e+02| 5.0e+02| 8.7e+02|
NGC7331         |CO6-5  | | 3.7e+02| 2.8e+02| 5.0e+02|
NGC7331         |CO7-6  | | 9.1e+01| 2.9e+01| 1.6e+02| 2.5e+02
NGC7331         |CO9-8  | | 2.4e+02| 4.7e+01| 5.6e+02| 9.2e+02
NGC7331         |CO11-10| | 2.7e+02| 7.3e+01| 4.7e+02| 9.2e+02
NGC7331         |CO12-11| | 3.0e+02| 7.0e+01| 5.6e+02| 1.0e+03
NGC7331         |NII    | | 1.2e+04| 1.1e+04| 1.2e+04|
UGC12150        |CI1-0  | | 6.1e+02| 3.6e+02| 8.4e+02| 1.4e+03
UGC12150        |CI2-1  | | 4.4e+02| 3.8e+02| 5.0e+02|
UGC12150        |CO5-4  | | 6.5e+02| 4.9e+02| 8.4e+02|
UGC12150        |CO6-5  | | 5.7e+02| 4.8e+02| 6.5e+02|
UGC12150        |CO7-6  | | 3.9e+02| 3.3e+02| 4.6e+02|
UGC12150        |CO8-7  | | 3.3e+02| 2.4e+02| 4.3e+02|
UGC12150        |CO9-8  | | 1.7e+02| 7.4e+01| 2.9e+02| 4.5e+02
UGC12150        |CO10-9 | | 1.8e+02| 8.8e+01| 2.7e+02| 4.3e+02
UGC12150        |CO11-10| | 6.6e+01| 1.4e+01| 1.6e+02| 2.6e+02
UGC12150        |CO13-12| | 8.6e+01| 2.6e+01| 1.7e+02| 2.7e+02
UGC12150        |NII    | | 1.3e+03| 1.2e+03| 1.3e+03|
IRAS 22491-1808 |CI2-1  | | 7.7e+01| 4.3e+01| 1.1e+02| 1.8e+02
IRAS 22491-1808 |CO5-4  | | 4.7e+02| 3.3e+02| 5.9e+02|
IRAS 22491-1808 |CO6-5  | | 2.6e+02| 1.8e+02| 3.2e+02|
IRAS 22491-1808 |CO7-6  | | 2.2e+02| 1.9e+02| 2.6e+02|
IRAS 22491-1808 |CO8-7  | | 3.0e+02| 2.5e+02| 3.3e+02|
IRAS 22491-1808 |CO9-8  | | 1.5e+02| 5.1e+01| 2.2e+02| 3.0e+02
IRAS 22491-1808 |CO10-9 | | 2.7e+02| 2.0e+02| 3.4e+02|
IRAS 22491-1808 |CO11-10| | 2.0e+02| 1.5e+02| 2.6e+02|
IRAS 22491-1808 |CO12-11| | 1.6e+02| 1.1e+02| 2.0e+02|
IRAS 22491-1808 |CO13-12| | 1.3e+02| 9.7e+01| 1.7e+02|
IRAS 22491-1808 |NII    | | 9.8e+01| 5.4e+01| 1.4e+02|
NGC7465         |CI1-0  | | 2.7e+02| 1.1e+02| 4.4e+02| 7.0e+02
NGC7465         |CI2-1  | | 2.4e+02| 1.6e+02| 3.1e+02|
NGC7465         |CO4-3  | | 3.4e+02| 1.5e+02| 5.1e+02| 9.0e+02
NGC7465         |CO5-4  | | 4.4e+02| 2.1e+02| 6.1e+02|
NGC7465         |CO6-5  | | 1.2e+02| 3.7e+01| 2.1e+02| 3.4e+02
NGC7465         |CO7-6  | | 6.1e+01| 1.9e+01| 1.2e+02| 2.3e+02
NGC7465         |CO8-7  | | 1.9e+02| 7.1e+01| 3.0e+02| 4.7e+02
NGC7465         |CO9-8  | | 1.5e+02| 3.8e+01| 2.8e+02| 4.7e+02
NGC7465         |CO10-9 | | 1.3e+02| 5.0e+01| 2.4e+02| 4.0e+02
NGC7465         |CO11-10| | 6.3e+01| 9.7e+00| 1.4e+02| 2.2e+02
NGC7465         |NII    | | 5.0e+02| 4.1e+02| 6.0e+02|
NGC7469         |CI1-0  | | 1.3e+03| 1.1e+03| 1.5e+03|
NGC7469         |CI2-1  | | 1.5e+03| 1.5e+03| 1.6e+03|
NGC7469         |CO4-3  | | 2.4e+03| 2.1e+03| 2.6e+03|
NGC7469         |CO5-4  | | 2.3e+03| 2.2e+03| 2.4e+03|
NGC7469         |CO6-5  | | 1.8e+03| 1.7e+03| 1.8e+03|
NGC7469         |CO7-6  | | 1.2e+03| 1.2e+03| 1.3e+03|
NGC7469         |CO8-7  | | 8.3e+02| 7.6e+02| 8.9e+02|
NGC7469         |CO9-8  | | 6.3e+02| 5.7e+02| 6.9e+02|
NGC7469         |CO10-9 | | 4.1e+02| 3.5e+02| 4.6e+02|
NGC7469         |CO11-10| | 3.0e+02| 2.5e+02| 3.5e+02|
NGC7469         |CO12-11| | 2.0e+02| 1.6e+02| 2.5e+02|
NGC7469         |CO13-12| | 2.0e+02| 1.3e+02| 2.6e+02|
NGC7469         |NII    | | 2.4e+03| 2.3e+03| 2.4e+03|
ESO148-IG002    |CI1-0  | | 1.6e+01| 2.0e+00| 3.8e+01| 8.2e+01
ESO148-IG002    |CI2-1  | | 1.9e+02| 1.6e+02| 2.2e+02|
ESO148-IG002    |CO5-4  | | 1.8e+02| 1.4e+02| 2.3e+02|
ESO148-IG002    |CO6-5  | | 2.6e+02| 2.2e+02| 3.0e+02|
ESO148-IG002    |CO7-6  | | 3.1e+02| 2.8e+02| 3.4e+02|
ESO148-IG002    |CO8-7  | | 3.4e+02| 3.0e+02| 3.8e+02|
ESO148-IG002    |CO9-8  | | 3.1e+02| 2.4e+02| 3.8e+02|
ESO148-IG002    |CO10-9 | | 2.6e+02| 2.1e+02| 3.0e+02|
ESO148-IG002    |CO11-10| | 2.1e+02| 1.7e+02| 2.6e+02|
ESO148-IG002    |CO12-11| | 1.4e+02| 1.0e+02| 1.7e+02|
ESO148-IG002    |CO13-12| | 1.8e+02| 1.4e+02| 2.2e+02|
ESO148-IG002    |NII    | | 3.7e+02| 3.3e+02| 4.1e+02|
IC5298          |CI1-0  | | 7.6e+02| 3.0e+02| 1.1e+03| 1.8e+03
IC5298          |CI2-1  | | 3.9e+02| 3.0e+02| 4.6e+02|
IC5298          |CO5-4  | | 7.7e+02| 5.4e+02| 1.0e+03|
IC5298          |CO6-5  | | 7.3e+02| 6.1e+02| 8.5e+02|
IC5298          |CO7-6  | | 3.9e+02| 3.1e+02| 4.6e+02|
IC5298          |CO8-7  | | 4.6e+02| 3.6e+02| 5.5e+02|
IC5298          |CO9-8  | | 3.0e+02| 2.0e+02| 4.1e+02|
IC5298          |CO10-9 | | 6.1e+01| 1.7e+01| 1.3e+02| 2.1e+02
IC5298          |CO11-10| | 8.5e+01| 2.8e+01| 1.5e+02| 2.8e+02
IC5298          |CO12-11| | 8.5e+01| 2.6e+01| 1.6e+02| 2.4e+02
IC5298          |CO13-12| | 8.1e+01| 2.1e+01| 1.6e+02| 2.5e+02
IC5298          |NII    | | 5.6e+02| 4.9e+02| 6.4e+02|
NGC7552         |CI1-0  | | 2.6e+03| 2.2e+03| 2.9e+03|
NGC7552         |CI2-1  | | 3.8e+03| 3.7e+03| 3.9e+03|
NGC7552         |CO4-3  | | 5.8e+03| 5.4e+03| 6.2e+03|
NGC7552         |CO5-4  | | 5.5e+03| 5.2e+03| 5.7e+03|
NGC7552         |CO6-5  | | 5.3e+03| 5.2e+03| 5.4e+03|
NGC7552         |CO7-6  | | 4.0e+03| 3.9e+03| 4.1e+03|
NGC7552         |CO8-7  | | 3.1e+03| 2.9e+03| 3.2e+03|
NGC7552         |CO9-8  | | 1.8e+03| 1.7e+03| 2.0e+03|
NGC7552         |CO10-9 | | 1.2e+03| 1.0e+03| 1.3e+03|
NGC7552         |CO11-10| | 9.1e+02| 8.0e+02| 1.0e+03|
NGC7552         |CO12-11| | 3.6e+02| 2.6e+02| 4.6e+02|
NGC7552         |CO13-12| | 2.5e+02| 9.9e+01| 4.1e+02| 6.2e+02
NGC7552         |NII    | | 7.1e+03| 7.0e+03| 7.2e+03|
NGC7591         |CI1-0  | | 5.2e+02| 2.0e+02| 8.2e+02| 1.2e+03
NGC7591         |CI2-1  | | 6.2e+02| 5.8e+02| 6.7e+02|
NGC7591         |CO4-3  | | 1.1e+03| 6.9e+02| 1.4e+03| 1.8e+03
NGC7591         |CO5-4  | | 2.7e+02| 1.0e+02| 5.3e+02| 7.9e+02
NGC7591         |CO6-5  | | 5.0e+02| 3.9e+02| 6.2e+02|
NGC7591         |CO7-6  | | 4.1e+02| 3.6e+02| 4.7e+02|
NGC7591         |CO8-7  | | 2.8e+02| 2.2e+02| 3.6e+02|
NGC7591         |CO9-8  | | 2.5e+02| 1.2e+02| 3.7e+02| 5.0e+02
NGC7591         |CO10-9 | | 2.6e+02| 1.6e+02| 3.5e+02|
NGC7591         |CO11-10| | 1.1e+02| 3.6e+01| 2.2e+02| 3.6e+02
NGC7591         |CO12-11| | 9.6e+01| 2.8e+01| 1.9e+02| 2.8e+02
NGC7591         |CO13-12| | 1.1e+02| 4.3e+01| 1.8e+02| 3.2e+02
NGC7591         |NII    | | 1.1e+03| 1.0e+03| 1.2e+03|
NGC7592         |CI1-0  | | 3.6e+02| 1.2e+02| 6.8e+02| 1.2e+03
NGC7592         |CI2-1  | | 4.1e+02| 3.3e+02| 4.7e+02|
NGC7592         |CO5-4  | | 5.1e+02| 2.4e+02| 7.3e+02|
NGC7592         |CO6-5  | | 5.6e+02| 4.3e+02| 6.6e+02|
NGC7592         |CO7-6  | | 3.2e+02| 2.4e+02| 4.0e+02|
NGC7592         |CO8-7  | | 3.1e+02| 2.0e+02| 4.1e+02|
NGC7592         |CO9-8  | | 4.2e+02| 2.8e+02| 5.7e+02|
NGC7592         |CO10-9 | | 1.2e+02| 4.2e+01| 1.9e+02| 4.2e+02
NGC7592         |CO11-10| | 7.7e+01| 2.1e+01| 1.6e+02| 2.9e+02
NGC7592         |CO13-12| | 9.7e+01| 2.5e+01| 1.9e+02| 3.0e+02
NGC7592         |NII    | | 9.8e+02| 8.9e+02| 1.1e+03|
NGC7582         |CI1-0  | | 2.2e+03| 1.9e+03| 2.4e+03|
NGC7582         |CI2-1  | | 2.7e+03| 2.7e+03| 2.8e+03|
NGC7582         |CO4-3  | | 4.2e+03| 3.9e+03| 4.5e+03|
NGC7582         |CO5-4  | | 4.0e+03| 3.8e+03| 4.2e+03|
NGC7582         |CO6-5  | | 3.4e+03| 3.3e+03| 3.5e+03|
NGC7582         |CO7-6  | | 2.3e+03| 2.3e+03| 2.4e+03|
NGC7582         |CO8-7  | | 1.8e+03| 1.6e+03| 1.9e+03|
NGC7582         |CO9-8  | | 1.4e+03| 1.3e+03| 1.6e+03|
NGC7582         |CO10-9 | | 8.6e+02| 7.7e+02| 9.6e+02|
NGC7582         |CO11-10| | 5.6e+02| 4.7e+02| 6.6e+02|
NGC7582         |CO12-11| | 2.1e+02| 1.2e+02| 2.9e+02| 4.1e+02
NGC7582         |CO13-12| | 2.5e+02| 9.3e+01| 4.1e+02| 6.3e+02
NGC7582         |NII    | | 4.0e+03| 3.9e+03| 4.2e+03|
IRAS 23230-6926 |CI2-1  | | 4.3e+01| 3.2e+01| 5.6e+01|
IRAS 23230-6926 |CO5-4  | | 2.6e+01| 9.5e+00| 4.9e+01| 8.0e+01
IRAS 23230-6926 |CO6-5  | | 4.2e+01| 2.1e+01| 6.1e+01| 8.1e+01
IRAS 23230-6926 |CO7-6  | | 5.7e+01| 4.5e+01| 7.2e+01|
IRAS 23230-6926 |CO8-7  | | 5.3e+01| 3.3e+01| 6.9e+01|
IRAS 23230-6926 |CO10-9 | | 1.2e+02| 7.9e+01| 1.7e+02|
IRAS 23230-6926 |CO11-10| | 7.1e+01| 3.8e+01| 1.0e+02| 1.5e+02
IRAS 23230-6926 |CO12-11| | 8.5e+01| 5.2e+01| 1.2e+02|
IRAS 23230-6926 |CO13-12| | 6.8e+01| 4.0e+01| 9.1e+01|
IRAS 23230-6926 |NII    | | 4.0e+01| 1.5e+01| 7.8e+01| 1.2e+02
NGC7674         |CI1-0  | | 1.1e+02| 2.0e+01| 2.0e+02| 3.7e+02
NGC7674         |CI2-1  | | 2.0e+02| 1.7e+02| 2.4e+02|
NGC7674         |CO5-4  | | 9.5e+01| 3.0e+01| 1.9e+02| 3.5e+02
NGC7674         |CO6-5  | | 1.1e+02| 5.6e+01| 1.6e+02| 2.4e+02
NGC7674         |CO7-6  | | 7.9e+01| 4.5e+01| 1.2e+02|
NGC7674         |CO8-7  | | 1.2e+02| 7.6e+01| 1.6e+02|
NGC7674         |CO9-8  | | 1.2e+02| 3.3e+01| 2.2e+02| 3.4e+02
NGC7674         |CO10-9 | | 8.6e+01| 2.2e+01| 1.5e+02| 2.6e+02
NGC7674         |CO11-10| | 8.1e+01| 2.1e+01| 1.5e+02| 2.4e+02
NGC7674         |CO12-11| | 1.8e+02| 1.1e+02| 2.5e+02|
NGC7674         |CO13-12| | 7.1e+01| 1.9e+01| 1.4e+02| 2.4e+02
NGC7674         |NII    | | 1.1e+03| 1.0e+03| 1.2e+03|
IRAS 23253-5415 |CI2-1  | | 7.0e+01| 4.1e+01| 9.9e+01|
IRAS 23253-5415 |CO5-4  | | 9.0e+01| 2.3e+01| 1.6e+02| 2.9e+02
IRAS 23253-5415 |CO6-5  | | 7.6e+01| 2.8e+01| 1.4e+02| 2.2e+02
IRAS 23253-5415 |CO7-6  | | 7.8e+01| 4.4e+01| 1.1e+02|
IRAS 23253-5415 |CO8-7  | | 6.4e+01| 3.9e+01| 9.0e+01|
IRAS 23253-5415 |CO10-9 | | 7.4e+01| 2.6e+01| 1.1e+02| 1.7e+02
IRAS 23253-5415 |CO11-10| | 4.2e+01| 1.5e+01| 7.4e+01| 1.0e+02
IRAS 23253-5415 |CO12-11| | 4.5e+01| 1.2e+01| 8.1e+01| 1.4e+02
IRAS 23253-5415 |CO13-12| | 5.0e+01| 1.8e+01| 8.7e+01| 1.3e+02
IRAS 23253-5415 |NII    | | 1.0e+02| 6.7e+01| 1.4e+02|
NGC7679a        |CI1-0  | | 4.8e+02| 1.5e+02| 8.0e+02| 1.2e+03
NGC7679a        |CI2-1  | | 2.8e+02| 2.0e+02| 3.6e+02|
NGC7679a        |CO4-3  | | 5.5e+02| 2.1e+02| 9.5e+02| 1.5e+03
NGC7679a        |CO5-4  | | 4.9e+02| 2.7e+02| 7.4e+02|
NGC7679a        |CO6-5  | | 6.8e+02| 5.7e+02| 7.9e+02|
NGC7679a        |CO7-6  | | 3.5e+02| 2.8e+02| 4.4e+02|
NGC7679a        |CO8-7  | | 1.5e+02| 5.6e+01| 2.4e+02| 3.7e+02
NGC7679a        |CO9-8  | | 4.6e+01| 4.9e+00| 1.6e+02| 2.8e+02
NGC7679a        |CO10-9 | | 2.0e+02| 9.9e+01| 2.9e+02| 4.4e+02
NGC7679a        |CO11-10| | 1.5e+02| 5.4e+01| 2.6e+02| 4.3e+02
NGC7679a        |CO12-11| | 2.0e+02| 1.0e+02| 2.8e+02|
NGC7679a        |CO13-12| | 1.2e+02| 3.4e+01| 2.2e+02| 3.7e+02
NGC7679a        |NII    | | 1.9e+03| 1.8e+03| 2.0e+03|
IRAS 23365+3604 |CI1-0  | | 4.2e+02| 1.8e+02| 6.8e+02| 1.1e+03
IRAS 23365+3604 |CI2-1  | | 2.4e+02| 1.9e+02| 2.8e+02|
IRAS 23365+3604 |CO5-4  | | 1.7e+02| 5.2e+01| 3.5e+02| 5.4e+02
IRAS 23365+3604 |CO6-5  | | 3.6e+02| 2.5e+02| 4.4e+02|
IRAS 23365+3604 |CO7-6  | | 3.5e+02| 3.0e+02| 4.1e+02|
IRAS 23365+3604 |CO8-7  | | 1.8e+02| 1.1e+02| 2.2e+02|
IRAS 23365+3604 |CO9-8  | | 1.5e+02| 4.9e+01| 2.5e+02| 3.8e+02
IRAS 23365+3604 |CO10-9 | | 2.9e+02| 2.2e+02| 3.6e+02|
IRAS 23365+3604 |CO11-10| | 1.4e+02| 6.5e+01| 1.9e+02| 2.8e+02
IRAS 23365+3604 |CO12-11| | 1.6e+02| 1.0e+02| 2.2e+02|
IRAS 23365+3604 |CO13-12| | 6.5e+01| 2.4e+01| 1.1e+02| 1.8e+02
IRAS 23365+3604 |NII    | | 1.9e+02| 1.4e+02| 2.5e+02|
NGC7771         |CI1-0  | | 1.0e+03| 8.8e+02| 1.2e+03|
NGC7771         |CI2-1  | | 1.1e+03| 1.1e+03| 1.2e+03|
NGC7771         |CO4-3  | | 1.6e+03| 1.5e+03| 1.8e+03|
NGC7771         |CO5-4  | | 1.6e+03| 1.5e+03| 1.7e+03|
NGC7771         |CO6-5  | | 1.3e+03| 1.3e+03| 1.4e+03|
NGC7771         |CO7-6  | | 7.3e+02| 6.9e+02| 7.8e+02|
NGC7771         |CO8-7  | | 5.3e+02| 4.6e+02| 6.0e+02|
NGC7771         |CO9-8  | | 3.6e+02| 2.9e+02| 4.2e+02|
NGC7771         |CO10-9 | | 1.5e+02| 9.9e+01| 2.0e+02| 2.5e+02
NGC7771         |CO11-10| | 2.0e+02| 1.5e+02| 2.6e+02|
NGC7771         |CO12-11| | 8.0e+01| 3.2e+01| 1.2e+02| 1.8e+02
NGC7771         |CO13-12| | 5.5e+01| 1.5e+01| 9.8e+01| 1.8e+02
NGC7771         |NII    |X| 5.6e+03| 5.5e+03| 5.7e+03|
Mrk331          |CI1-0  | | 8.9e+02| 6.9e+02| 1.0e+03|
Mrk331          |CI2-1  | | 7.3e+02| 7.0e+02| 7.7e+02|
Mrk331          |CO5-4  | | 1.1e+03| 1.0e+03| 1.2e+03|
Mrk331          |CO6-5  | | 1.0e+03| 9.6e+02| 1.0e+03|
Mrk331          |CO7-6  | | 6.6e+02| 6.3e+02| 7.0e+02|
Mrk331          |CO8-7  | | 4.6e+02| 4.2e+02| 5.1e+02|
Mrk331          |CO9-8  | | 4.7e+02| 4.2e+02| 5.2e+02|
Mrk331          |CO10-9 | | 2.4e+02| 1.9e+02| 2.8e+02|
Mrk331          |CO11-10| | 2.0e+02| 1.6e+02| 2.5e+02|
Mrk331          |CO12-11| | 1.3e+02| 1.0e+02| 1.6e+02|
Mrk331          |CO13-12| | 1.3e+02| 8.6e+01| 1.6e+02|
Mrk331          |NII    |X| 2.2e+03| 2.1e+03| 2.2e+03|
