ID                           LIR4-120[Lsun]   DL[Mpc]                   Redshift
NGC0023                     |  10.9       |     68                 |     0.015231
NGC0034                     |  11.2       |     85                 |    0.019617
MCG-02-01-051               |  11.2       |     120                |    0.027103
IC10                        |  7.5        |     1                  |    -0.001161
IRAS00188-0856              |  12.2       |     591                |    0.12842
ESO350-IG038                |  10.8       |     87                 |    0.020598
NGC205                      |  6.1        |     1                  |    -0.000804
IRAS00397-1312              |  12.6       |     1285               |    0.261717
NGC0232a                    |  11.2       |     95                 |    0.022639
NGC253                      |  10.3       |     3                  |    0.000811
IZw1                        |  11.4       |     272                |    0.0589
MCG+12-02-001               |  11.2       |     72                 |    0.015698
NGC0317B                    |  11.0       |     80                 |    0.018109
IRAS01003-2238              |  11.9       |     539                |    0.117835
3C31                        |             |     75                 |    0.017005
IC1623                      |  11.4       |     86                 |    0.020067
MCG-03-04-014               |  11.4       |     152                |    0.035144
ESO244-G012                 |  11.1       |     95                 |    0.022903
CGCG436-030                 |  11.5       |     138                |    0.031229
ESO353-G020                 |  10.8       |     66                 |    0.015921
IIIZw035                    |             |     120                |    0.027436
NGC0695                     |  11.4       |     143                |    0.032472
Mrk1014                     |  12.3       |     763                |    0.16311
NGC0828                     |  11.1       |     80                 |    0.017926
NGC0877                     |             |     57                 |    0.013052
NGC891                      |  10.2       |     10                 |    0.001761
UGC01845                    |  10.9       |     70                 |    0.015607
NGC0958                     |  10.9       |     82                 |    0.01914
0235+164                    |             |     4278               |    0.94
NGC1068                     |  10.9       |     16                 |    0.003793
NGC1056                     |  9.7        |     24                 |    0.005154
UGC02238                    |  11.1       |     93                 |    0.021883
NGC1097                     |  10.4       |     16                 |    0.00424
UGC02369                    |  11.4       |     142                |    0.031202
NGC1222                     |  10.4       |     35                 |    0.008079
UGC02608                    |  11.1       |     104                |    0.023343
NGC1266                     |  10.2       |     31                 |    0.007238
IRAS03158+4227              |  12.4       |     623                |    0.13443
3C84                        |  10.8       |     78                 |    0.017559
NGC1365-SW                  |  10.8       |     21                 |    0.005457
NGC1365-NE                  |  10.8       |     21                 |    0.005457
NGC1377                     |  9.7        |     24                 |    0.005977
NGC1482                     |  10.5       |     25                 |    0.006391
IRAS03521+0028              |  12.3       |     709                |    0.15191
UGC02982                    |  10.9       |     77                 |    0.017696
ESO420-G013                 |  10.7       |     49                 |    0.011908
NGC1572                     |  11.0       |     86                 |    0.020384
IRAS04271+3849              |  10.9       |     86                 |    0.018813
NGC1614                     |  11.3       |     68                 |    0.015938
UGC03094                    |  11.1       |     108                |    0.02471
MCG-05-12-006               |  10.9       |     78                 |    0.018753
IRASF05189-2524             |  11.8       |     185                |    0.042563
IRAS05223+1908              |             |     130                |    0.029577
MCG+08-11-002               |  11.2       |     86                 |    0.019157
NGC1961                     |  10.7       |     61                 |    0.013122
UGC03351                    |  11.1       |     67                 |    0.01486
IRAS05442+1732              |  11.0       |     81                 |    0.01862
IRAS06035-7102              |  12.0       |     353                |    0.079465
UGC03410a                   |  10.8       |     61                 |    0.013079
NGC2146-NW                  |  10.8       |     17                 |    0.002979
NGC2146-nuc                 |  10.8       |     17                 |    0.002979
NGC2146-SE                  |  10.8       |     17                 |    0.002979
IRAS06206-6315              |  12.0       |     411                |    0.092441
ESO255-IG007                |             |     166                |    0.03879
UGC03608                    |  11.1       |     97                 |    0.021351
NGC2342b                    |  10.8       |     77                 |    0.017599
NGC2342a                    |  10.8       |     77                 |    0.017599
NGC2369                     |  10.8       |     43                 |    0.010807
NGC2388a                    |  11.0       |     62                 |    0.01379
MCG+02-20-003               |  10.8       |     72                 |    0.016255
IRAS07598+6508              |  12.1       |     693                |    0.1483
B20827+24                   |             |     5818               |    0.9414
IRAS08311-2459              |  12.2       |     451                |    0.100449
He2-10                      |  9.6        |     10                 |    0.002912
IRAS08355-4944              |             |     110                |    0.025898
NGC2623                     |  11.4       |     81                 |    0.018509
IRAS08572+3915              |  11.8       |     261                |    0.05835
IRAS09022-3615              |  12.0       |     262                |    0.059641
NGC2764                     |  10.0       |     40                 |    0.009026
NGC2798                     |  10.4       |     28                 |    0.005757
UGC05101                    |  11.8       |     176                |    0.039367
NGC2976_00                  |             |     4                  |    1e-05
M81                         |  9.2        |     4                  |    -0.000113
M82                         |  10.4       |     4                  |    0.000677
NGC3077                     |  7.7        |     1                  |    4.7e-05
NGC3110a                    |  11.0       |     73                 |    0.016858
3C236                       |             |     451                |    0.1005
NGC3221                     |  10.7       |     61                 |    0.013709
NGC3227                     |  9.7        |     18                 |    0.003859
NGC3256                     |  11.3       |     38                 |    0.009354
IRAS10378+1109              |  12.1       |     631                |    0.136274
ESO264-G036                 |  10.9       |     89                 |    0.021065
NGC3351                     |  9.7        |     13                 |    0.002595
ESO264-G057                 |  10.7       |     72                 |    0.017199
IRASF10565+2448             |  11.8       |     192                |    0.0431
NGC3521                     |  10.1       |     12                 |    0.002672
IRAS11095-0238              |  12.0       |     482                |    0.106634
NGC3627                     |  10.2       |     12                 |    0.002425
NGC3665                     |  9.7        |     32                 |    0.006901
Arp299-B                    |  11.6       |     49                 |    0.0103
Arp299-C                    |  11.6       |     49                 |    0.0103
Arp299-A                    |  11.6       |     49                 |    0.0103
PG1126-041                  |             |     266                |    0.06196
ESO320-G030                 |  11.0       |     45                 |    0.010781
NGC3982                     |  9.8        |     21                 |    0.003699
NGC4038                     |             |     23                 |    0.005477
NGC4038overlap              |             |     23                 |    0.005477
NGC4051                     |  9.5        |     14                 |    0.002336
IRAS12071-0444              |  12.1       |     591                |    0.128355
NGC4151                     |             |     18                 |    0.003319
NGC4194                     |  10.7       |     39                 |    0.008342
IRAS12116-5615              |  11.3       |     115                |    0.027102
NGC4254                     |  10.8       |     36                 |    0.008029
NGC4321                     |  10.4       |     25                 |    0.00524
NGC4388                     |  10.4       |     38                 |    0.008419
NGC4459                     |  9.1        |     19                 |    0.003976
NGC4526                     |  9.1        |     10                 |    0.002058
NGC4536                     |  10.5       |     27                 |    0.006031
NGC4569                     |  7.5        |     1                  |    -0.000784
TOL1238-364                 |  10.4       |     46                 |    0.010924
NGC4631                     |  10.4       |     12                 |    0.002021
NGC4710                     |  9.6        |     18                 |    0.003676
NGC4736                     |  9.9        |     8                  |    0.001027
Mrk231                      |  12.2       |     188                |    0.04217
NGC4826                     |  9.7        |     9                  |    0.001361
MCG-02-33-098               |  10.7       |     69                 |    0.015921
ESO507-G070                 |  11.2       |     91                 |    0.021702
NGC5010                     |  10.6       |     43                 |    0.009924
IRAS13120-5453              |  12.0       |     132                |    0.030761
NGC5055                     |  10.1       |     11                 |    0.001614
Arp193                      |  11.4       |     105                |    0.023299
NGC5104                     |  10.9       |     82                 |    0.018606
MCG-03-34-064               |             |     74                 |    0.016541
CenA                        |  9.7        |     4                  |    0.001825
NGC5135                     |  11.0       |     58                 |    0.013693
ESO173-G015                 |  11.2       |     39                 |    0.009735
NGC5194                     |  10.4       |     11                 |    0.001544
IC4280                      |  10.7       |     70                 |    0.016308
M83                         |  10.4       |     7                  |    0.001711
Mrk273                      |  12.0       |     168                |    0.03778
4C12.50                     |  12.0       |     561                |    0.12174
UGC08739                    |  10.8       |     76                 |    0.016785
ESO221-IG010                |  10.5       |     39                 |    0.010337
Mrk463                      |  11.2       |     226                |    0.050355
M101_02                     |  10.1       |     8                  |    0.000804
OQ208                       |             |     348                |    0.076576
NGC5653                     |  10.8       |     55                 |    0.011881
IRAS14348-1447              |  12.1       |     371                |    0.083
NGC5713                     |  10.5       |     29                 |    0.006334
IRAS14378-3651              |  11.9       |     303                |    0.067637
Mrk478                      |  11.1       |     358                |    0.079055
NGC5734a                    |  10.7       |     59                 |    0.013746
3C305                       |             |     187                |    0.041639
VV340a                      |             |     145                |    0.033669
IC4518ABa                   |             |     68                 |    0.015728
NGC5866                     |  9.4        |     14                 |    0.002518
CGCG049-057                 |  11.1       |     59                 |    0.012999
3C315                       |             |     498                |    0.1083
VV705                       |             |     181                |    0.040191
ESO099-G004                 |  11.4       |     125                |    0.029284
IRAS15250+3609              |  11.8       |     248                |    0.055155
NGC5936                     |  10.8       |     61                 |    0.013356
Arp220                      |  12.0       |     81                 |    0.018126
NGC5990                     |  10.7       |     57                 |    0.012806
IRAS15462-0450              |  12.0       |     456                |    0.099792
3C326                       |             |     407                |    0.0895
PKS1549-79                  |             |     690                |    0.1522
NGC6052                     |  10.8       |     71                 |    0.015808
IRAS16090-0139              |  12.3       |     618                |    0.13358
PG1613+658                  |  11.5       |     600                |    0.129
CGCG052-037                 |  11.1       |     109                |    0.02449
NGC6156                     |  10.8       |     45                 |    0.010885
ESO069-IG006                |  11.7       |     203                |    0.046439
IRASF16399-0937             |  11.3       |     118                |    0.027012
NGC6240                     |  11.6       |     108                |    0.02448
IRASF16516-0948             |  11.0       |     100                |    0.022706
NGC6286b                    |  11.1       |     85                 |    0.018349
NGC6286a                    |  11.1       |     85                 |    0.018349
IRASF17138-1017             |  11.1       |     76                 |    0.017335
IRASF17208-0014             |  12.2       |     190                |    0.04281
ESO138-G027                 |  11.1       |     88                 |    0.020781
UGC11041                    |  10.8       |     74                 |    0.016281
IRAS17578-0400              |  11.2       |     62                 |    0.014043
NGC6621                     |  11.0       |     92                 |    0.020652
IC4687                      |  11.1       |     73                 |    0.017345
IRASF18293-3413             |  11.5       |     78                 |    0.018176
IC4734                      |  11.0       |     67                 |    0.015611
NGC6701                     |  10.9       |     62                 |    0.013226
IRAS19254-7245              |  11.8       |     270                |    0.061709
IRAS19297-0406              |  12.2       |     387                |    0.08573
ESO339-G011                 |  10.8       |     82                 |    0.0192
3C405                       |             |     252                |    0.056075
IRAS20087-0308              |  12.2       |     480                |    0.10567
IRAS20100-4156              |  12.4       |     595                |    0.129583
MCG+04-48-002a              |  10.9       |     65                 |    0.0139
NGC6926                     |  11.0       |     87                 |    0.019613
NGC6946                     |  9.8        |     5                  |    0.000133
NGC6946_05                  |  9.8        |     5                  |    0.000133
IRAS20414-1651              |  12.0       |     392                |    0.087084
3C424                       |             |     586                |    0.126988
IC5063                      |  10.2       |     46                 |    0.011348
CGCG448-020                 |  11.7       |     161                |    0.036098
ESO286-IG019                |  11.8       |     185                |    0.042996
ESO286-G035                 |  10.8       |     73                 |    0.017361
3C433                       |             |     465                |    0.1016
NGC7130                     |  11.1       |     69                 |    0.016151
NGC7172                     |  10.2       |     36                 |    0.008683
ESO467-G027                 |  10.8       |     74                 |    0.017401
IC5179                      |  10.9       |     48                 |    0.011415
NGC7331                     |  10.3       |     15                 |    0.002722
UGC12150                    |  11.1       |     96                 |    0.021391
IRAS22491-1808              |  11.9       |     345                |    0.07776
NGC7465                     |  9.7        |     30                 |    0.006538
NGC7469                     |  11.3       |     72                 |    0.016317
ESO148-IG002                |  11.8       |     193                |    0.044601
IC5298                      |  11.3       |     122                |    0.027422
NGC7552                     |  10.7       |     21                 |    0.005365
NGC7591                     |  10.8       |     72                 |    0.016531
NGC7592                     |  11.1       |     106                |    0.024444
NGC7582                     |  10.5       |     21                 |    0.005254
IRAS23230-6926              |  12.1       |     482                |    0.10659
NGC7674                     |  11.2       |     130                |    0.028924
IRAS23253-5415              |  12.1       |     595                |    0.13004
NGC7679                     |  10.8       |     75                 |    0.017139
IRAS23365+3604              |  12.0       |     290                |    0.06448
NGC7771                     |  11.1       |     63                 |    0.014267
Mrk331                      |  11.2       |     81                 |    0.018483
