#
#   VizieR Astronomical Server vizier.cfa.harvard.edu
#    Date: 2020-03-23T11:44:54 [V1.99+ (14-Oct-2013)]
#   In case of problem, please report to:	cds-question@unistra.fr
#
#
#Coosys	J2000:	eq_FK5 J2000
#INFO	votable-version=1.99+ (14-Oct-2013)	
#INFO	-ref=VIZ5e789c6310448	
#INFO	-out.max=unlimited	
#INFO	queryParameters=18	
#-oc.form=dec
#-out.max=unlimited
#-out.all=2
#-order=I
#-out.src=J/ApJ/829/93/table3
#-nav=cat:J/ApJ/829/93&tab:{J/ApJ/829/93/table3}&key:source=J/ApJ/829/93/table3&HTTPPRM:&&-ref=VIZ5e789c6310448&-out.max=unlimited&-out.form=HTML Table&-oc.form=sexa&-order=I&-out=ID&-out=Jup&-out=RFlux&-out=sigmam&-out=sigmac&-out=x_RFlux&-out=dv&-out=Omegab&-out=Flux&-out=e_Flux&-out=r_RFlux&-file=.&-meta.ucd=2&-meta=1&-meta.foot=1&-usenav=1&-bmark=POST&-out.src=J/ApJ/829/93/table3
#-source=J/ApJ/829/93/table3
#-out=ID
#-out=Jup
#-out=RFlux
#-out=sigmam
#-out=sigmac
#-out=x_RFlux
#-out=dv
#-out=Omegab
#-out=Flux
#-out=e_Flux
#-out=r_RFlux
#

#RESOURCE=yCat_18290093
#Name: J/ApJ/829/93
#Title: CO, [CI] and [NII] lines from Herschel spectra (Kamenetzky+, 2016)
#Table	J_ApJ_829_93_table3:
#Name: J/ApJ/829/93/table3
#Title: CO J=1-0 to J=3-2 line fluxes
#Column	ID	(a19)	Galaxy identifier	[ucd=meta.id;meta.main]
#Column	Jup	(I1)	[1/7] Upper J level	[ucd=phys.atmol.qn]
#Column	RFlux	(E9.2)	[0/28600] Reported line flux	[ucd=phot.flux]
#Column	sigmam	(E9.2)	[0/3400] Measurement error in RFlux (1)	[ucd=stat.error]
#Column	sigmac	(E9.2)	[0/2950] Calibration error in RFlux (1)	[ucd=stat.error]
#Column	x_RFlux	(A5)	Units of RFlux (2)	[ucd=meta.unit]
#Column	dv	(I3)	[11/580]? Line velocity Full-Width at Half-Maximum [NULL integer written as an empty string]	[ucd=spect.line.width]
#Column	Omegab	(I2)	[8/55]? Beam size Full-Width at Half-Maximum [NULL integer written as an empty string]	[ucd=phys.angSize]
#Column	Flux	(E9.2)	[0/89300]? This analysis line flux (3)	[ucd=phot.flux.density;spect.line]
#Column	e_Flux	(E9.2)	[0.3/26800]? Total uncertainty in Flux (3)	[ucd=stat.error;phot.flux]
#Column	r_RFlux	(I2)	Reference for RFlux (see refs.dat file)	[ucd=meta.ref;pos.frame]
ID|Jup|RFlux|sigmam|sigmac|x_RFlux|dv|Omegab|Flux|e_Flux|r_RFlux
 | | | | | |km/s|arcsec|Jy.km/s|Jy.km/s|
-------------------|-|---------|---------|---------|-----|---|--|---------|---------|--
NGC0023            |1| 1.69e+01| 0.00e+00| 4.22e+00|Kkms |141|24| 1.39e+02| 3.47e+01| 1
NGC0023            |1| 6.00e+00| 0.00e+00| 1.20e+00|Kkms |374|55| 1.70e+02| 3.40e+01| 2
NGC0023            |1| 8.90e+00| 0.00e+00| 2.23e+00|Kkms |190|45| 1.84e+02| 4.61e+01| 1
NGC0023            |1| 1.80e+01| 0.00e+00| 1.30e+00|Kkms |   |33| 2.34e+02| 1.69e+01| 3
NGC0023            |1| 3.40e+01| 3.84e-01| 6.81e+00|Kkms |   |22| 2.47e+02| 4.96e+01| 4
NGC0023            |2| 1.88e+01| 0.00e+00| 4.70e+00|Kkms |129|12| 2.36e+02| 5.89e+01| 1
NGC0023            |2| 7.40e+00| 0.00e+00| 1.85e+00|Kkms |210|24| 2.43e+02| 6.08e+01| 1
NGC0023            |3| 1.53e+01| 1.27e+00| 2.30e+00|Kkms |257|22| 1.00e+03| 1.72e+02| 5
NGC34              |1| 1.70e+01| 0.00e+00| 4.25e+00|Kkms |149|24| 1.15e+02| 2.88e+01| 1
NGC34              |1| 4.49e+00| 3.10e-01| 4.49e-01|Kkms |295|55| 1.32e+02| 1.60e+01| 6
NGC34              |1| 6.70e+00| 0.00e+00| 1.68e+00|Kkms |274|45| 1.38e+02| 3.46e+01| 1
NGC34              |1| 1.48e+02| 1.35e+01| 2.97e+01|Jykms|   |45| 1.48e+02| 3.24e+01| 7
NGC34              |2| 4.30e+00| 0.00e+00| 1.07e+00|Kkms |271|24| 1.17e+02| 2.92e+01| 1
NGC34              |2| 5.65e+01| 0.00e+00| 1.41e+01|Kkms |172|12| 4.72e+02| 1.18e+02| 1
NGC34              |3| 7.70e+00| 1.76e+00| 1.16e+00|Kkms |168|22| 4.05e+02| 1.11e+02| 5
MCG-02-01-051      |1| 2.29e+00| 2.52e-01| 3.44e-01|Kkms |266|55| 6.31e+01| 1.17e+01| 8
MCG-02-01-051      |2| 5.32e+00| 4.47e-01| 7.99e-01|Kkms |247|32| 2.41e+02| 4.14e+01| 5
IC10-B11-1         |1| 8.10e+00| 0.00e+00| 8.10e-01|Kkms | 11|55| 2.04e+02| 2.04e+01| 9
IC10-B11-1         |2| 1.33e+01| 7.30e-01| 1.99e+00|Kkms | 36|32| 8.53e+02| 1.36e+02| 5
IC10-B11-1         |2| 2.23e+01| 2.00e-01| 2.23e+00|Kkms |   |30| 1.38e+03| 1.38e+02|10
IC10-B11-1         |3| 7.10e+00| 3.00e-01| 2.13e+00|Kkms | 14|22| 7.56e+02| 2.29e+02|11
IC10-B11-1         |3| 1.27e+01| 7.00e-01| 1.27e+00|Kkms |   |21| 1.35e+03| 1.54e+02|10
IC10-B11-1         |4| 1.04e+01| 1.20e+00| 1.04e+00|Kkms |   |14| 1.40e+03| 2.14e+02|10
IC10-B11-1         |6| 3.10e+00| 5.00e+00| 3.10e-01|Kkms |   |10| 7.23e+02| 1.17e+03|10
IC10-B11-1         |7| 3.60e+00| 8.00e-01| 3.60e-01|Kkms |   | 8| 9.94e+02| 2.42e+02|10
NGC0232a           |1| 8.90e+00| 0.00e+00| 1.78e+00|Kkms |   |44| 1.75e+02| 3.50e+01|12
NGC0232a           |1| 2.10e+02| 5.70e+00| 4.20e+01|Jykms|   |45| 2.09e+02| 4.21e+01| 7
NGC0232a           |1| 1.11e+01| 3.00e-01| 1.11e+00|Kkms |358|45| 2.27e+02| 2.35e+01|13
NGC0232a           |1| 1.15e+01| 0.00e+00| 2.88e+00|Kkms |433|45| 2.36e+02| 5.89e+01| 1
NGC0232a           |1| 3.82e+01| 0.00e+00| 9.55e+00|Kkms |162|24| 2.53e+02| 6.32e+01| 1
NGC0232a           |2| 5.13e+01| 0.00e+00| 1.28e+01|Kkms |178|12| 4.03e+02| 1.01e+02| 1
NGC0232a           |2| 1.58e+01| 4.00e-01| 1.58e+00|Kkms |309|24| 4.18e+02| 4.31e+01|13
NGC0232a           |2| 1.78e+01| 0.00e+00| 4.45e+00|Kkms | 88|24| 4.71e+02| 1.18e+02| 1
NGC0232a           |2| 3.24e+02| 8.20e+00| 6.48e+01|Jykms|   |  |         |         | 7
NGC253             |1| 9.20e+02| 0.00e+00| 8.28e+01|Kkms |   |23| 7.06e+03| 6.36e+02|14
NGC253             |1| 1.08e+04| 1.35e+02| 1.08e+03|Jykms|220|45| 1.06e+04| 1.07e+03|15
NGC253             |1| 8.24e+03| 0.00e+00| 1.65e+03|Jykms|   |  |         |         | 7
NGC253             |2| 2.86e+04| 1.80e+02| 2.86e+03|Jykms|   |33| 3.22e+04| 3.23e+03|16
NGC253             |2| 1.06e+03| 0.00e+00| 1.17e+02|Kkms |   |23| 3.26e+04| 3.59e+03|14
NGC253             |3| 9.98e+02| 0.00e+00| 1.40e+02|Kkms |   |23| 6.90e+04| 9.65e+03|14
IZw1               |1| 0.00e+00| 5.90e-01| 0.00e+00|Kkms |   |55| 0.00e+00| 1.53e+01| 6
IZw1               |1| 7.00e+00| 0.00e+00| 1.40e+00|Kkms |410|22| 3.57e+01| 7.14e+00|17
IZw1               |1| 3.40e+01| 7.00e+00| 5.10e+00|Jykms|   |  |         |         |18
IZw1               |2| 1.14e+02| 2.30e+01| 1.71e+01|Jykms|   |  |         |         |18
IZw1               |3| 3.56e+02| 1.03e+02| 5.34e+01|Jykms|   |  |         |         |18
IZw1               |6| 4.30e+02| 1.55e+02| 1.08e+02|Jykms|   | 8| 5.99e+02| 2.63e+02|18
MCG+12-02-001      |1| 4.38e+01| 4.68e-01| 8.76e+00|Kkms |   |22| 2.87e+02| 5.76e+01| 4
MCG+12-02-001      |2| 2.63e+01| 5.99e-01| 3.95e+00|Kkms |231|32| 1.24e+03| 1.88e+02| 5
MCG+12-02-001      |3| 2.87e+01| 1.14e+00| 4.31e+00|Kkms |183|22| 1.70e+03| 2.63e+02| 5
NGC0317B           |1| 4.21e+00| 2.34e-01| 6.32e-01|Kkms |275|55| 1.24e+02| 1.98e+01| 8
NGC0317B           |2| 1.94e+01| 6.95e-01| 2.90e+00|Kkms |386|32| 8.78e+02| 1.35e+02| 5
NGC0317B           |3| 1.19e+01| 6.68e-01| 1.79e+00|Kkms |255|22| 6.33e+02| 1.01e+02| 5
3C 31              |1| 2.70e+01| 2.00e+00| 4.05e+00|Jykms|450|55| 2.55e+01| 4.26e+00|19
IC1623             |1| 1.74e+01| 5.71e-01| 1.74e+00|Kkms |   |34| 2.30e+02| 2.43e+01|20
IC1623             |1| 1.41e+01| 0.00e+00| 2.82e+00|Kkms |237|55| 3.98e+02| 7.96e+01| 2
IC1623             |1| 6.91e+02| 1.38e+02| 1.04e+02|Jykms|   |  |         |         |18
IC1623             |1| 2.91e+02| 4.48e+01| 5.82e+01|Jykms|   |  |         |         | 7
IC1623             |2| 3.52e+01| 9.21e-01| 5.29e+00|Kkms |279|32| 1.70e+03| 2.59e+02| 5
IC1623             |3| 4.51e+01| 1.76e+00| 6.76e+00|Kkms |297|22| 2.95e+03| 4.57e+02| 5
IC1623             |3| 1.08e+02| 0.00e+00| 2.16e+01|Kkms |301|14| 4.25e+03| 8.49e+02|21
IC1623             |3| 3.32e+03| 6.60e+02| 4.99e+02|Jykms|   |  |         |         |18
MCG-03-04-014      |1| 4.90e+00| 0.00e+00| 9.80e-01|Kkms |   |44| 9.29e+01| 1.86e+01|12
MCG-03-04-014      |1| 1.20e+02| 0.00e+00| 2.40e+01|Jykms|   |45| 1.19e+02| 2.39e+01| 7
MCG-03-04-014      |1| 1.78e+02| 3.60e+01| 2.67e+01|Jykms|   |  |         |         |18
MCG-03-04-014      |2| 6.69e+00| 2.46e-01| 1.00e+00|Kkms |280|32| 2.85e+02| 4.40e+01| 5
MCG-03-04-014      |3| 4.79e+00| 6.43e-01| 7.18e-01|Kkms |154|22| 2.39e+02| 4.82e+01| 5
MCG-03-04-014      |3| 1.53e+01| 0.00e+00| 3.06e+00|Kkms |230|14| 3.59e+02| 7.17e+01|21
MCG-03-04-014      |3| 5.07e+02| 1.00e+02| 7.60e+01|Jykms|   |  |         |         |18
ESO244-G012        |1| 4.40e+00| 0.00e+00| 8.80e-01|Kkms |   |44| 8.63e+01| 1.73e+01|12
ESO244-G012        |1| 1.08e+02| 0.00e+00| 2.16e+01|Jykms|   |45| 1.06e+02| 2.13e+01| 7
ESO244-G012        |1| 6.30e+00| 0.00e+00| 1.57e+00|Kkms |275|45| 1.28e+02| 3.20e+01| 1
ESO244-G012        |2| 1.43e+01| 0.00e+00| 3.58e+00|Kkms |201|24| 4.54e+02| 1.14e+02| 1
CGCG436-030        |2| 6.20e+00| 4.06e-01| 9.30e-01|Kkms |216|32| 2.69e+02| 4.40e+01| 5
CGCG436-030        |3| 9.84e+00| 6.66e-01| 1.48e+00|Kkms |180|22| 5.09e+02| 8.38e+01| 5
IRASF01417+1651    |1| 1.80e+00| 0.00e+00| 3.60e-01|Kkms |164|55| 5.24e+01| 1.05e+01| 2
IRASF01417+1651    |1| 1.25e+01| 4.20e-01| 2.50e+00|Kkms |   |22| 6.74e+01| 1.37e+01| 4
IRASF01417+1651    |1| 7.50e+01| 1.50e+01| 1.12e+01|Jykms|   |  |         |         |18
IRASF01417+1651    |2| 6.42e+00| 4.06e-01| 9.63e-01|Kkms |240|32| 2.76e+02| 4.49e+01| 5
IRASF01417+1651    |3| 4.40e+00| 6.00e-01| 1.32e+00|Kkms |141|22| 2.13e+02| 7.03e+01|11
IRASF01417+1651    |3| 1.85e+01| 0.00e+00| 3.70e+00|Kkms |262|14| 3.90e+02| 7.81e+01|21
IRASF01417+1651    |3| 4.17e+02| 8.30e+01| 6.25e+01|Jykms|   |  |         |         |18
NGC0695            |1| 2.73e+01| 0.00e+00| 5.46e+00|Jykms|   |21| 3.59e+01| 7.18e+00| 7
NGC0695            |1| 6.00e+00| 0.00e+00| 1.20e+00|Kkms |300|55| 1.67e+02| 3.34e+01| 2
NGC0695            |2| 1.50e+01| 6.35e-01| 2.25e+00|Kkms |201|32| 6.68e+02| 1.04e+02| 5
NGC0695            |3| 1.35e+01| 9.26e-01| 2.02e+00|Kkms |184|22| 7.47e+02| 1.23e+02| 5
Mrk 1014           |1| 1.80e+00| 0.00e+00| 6.30e-01|Kkms |200|22| 7.02e+00| 2.46e+00|17
NGC0828            |1| 1.23e+01| 0.00e+00| 2.46e+00|Kkms |300|55| 3.57e+02| 7.14e+01| 2
NGC0828            |1| 3.78e+02| 0.00e+00| 7.56e+01|Jykms|   |21| 4.90e+02| 9.81e+01| 7
NGC0828            |1| 5.00e+01| 2.00e+00| 5.00e+00|Kkms |   |33| 6.11e+02| 6.58e+01|20
NGC0828            |1| 4.08e+02| 3.30e+01| 6.12e+01|Jykms|   |  |         |         |18
NGC0828            |2| 1.24e+03| 2.48e+02| 1.86e+02|Jykms|   |  |         |         |18
NGC0828            |3| 2.56e+03| 5.15e+02| 3.84e+02|Jykms|   |  |         |         |18
NGC0877a           |1| 1.22e+01| 0.00e+00| 3.05e+00|Kkms |143|24| 1.55e+02| 3.88e+01| 1
NGC0877a           |1| 9.10e+00| 0.00e+00| 1.82e+00|Kkms |200|55| 2.25e+02| 4.50e+01| 2
NGC0877a           |1| 1.16e+01| 0.00e+00| 2.90e+00|Kkms |342|45| 2.37e+02| 5.91e+01| 1
NGC0877a           |2| 1.04e+01| 0.00e+00| 2.60e+00|Kkms |213|24| 5.30e+02| 1.32e+02| 1
NGC0877a           |2| 1.29e+01| 0.00e+00| 3.23e+00|Kkms |132|12| 5.33e+02| 1.33e+02| 1
NGC891-1           |1| 3.73e+01| 9.20e-01| 5.59e+00|Kkms |172|55| 9.79e+02| 1.49e+02| 8
NGC891-1           |1| 4.94e+02| 0.00e+00| 9.89e+01|Jykms|   |  |         |         | 7
NGC891-1           |2| 7.24e+01| 6.68e-01| 1.09e+01|Kkms |154|32| 4.25e+03| 6.39e+02| 5
NGC891-1           |2| 3.82e+02| 2.66e+01| 7.63e+01|Jykms|   |  |         |         | 7
NGC891-1           |3| 1.10e+01| 3.00e-01| 1.10e+00|Kkms |   |21| 9.76e+02| 1.01e+02|10
NGC891-1           |3| 1.73e+01| 1.00e+00| 5.19e+00|Kkms | 59|22| 1.54e+03| 4.71e+02|11
NGC891-1           |3| 4.86e+01| 2.15e+00| 7.29e+00|Kkms |118|22| 4.33e+03| 6.77e+02| 5
UGC01845           |1| 3.95e+01| 3.72e-01| 7.90e+00|Kkms |   |22| 2.21e+02| 4.43e+01| 4
UGC01845           |2| 2.20e+01| 7.53e-01| 3.30e+00|Kkms |387|32| 9.78e+02| 1.50e+02| 5
UGC01845           |3| 1.89e+01| 5.22e-01| 2.84e+00|Kkms |341|22| 9.55e+02| 1.46e+02| 5
NGC0958            |1| 7.40e+00| 0.00e+00| 1.48e+00|Kkms |239|55| 1.93e+02| 3.86e+01| 2
NGC1068            |1| 2.31e+03| 2.44e+02| 2.31e+02|Jykms|280|45| 2.25e+03| 3.27e+02|15
NGC1068            |1| 1.90e+03| 0.00e+00| 3.81e+02|Jykms|   |21| 4.18e+03| 8.36e+02| 7
NGC1068            |1| 2.83e+03| 4.24e+02| 4.24e+02|Jykms|   |  |         |         |18
NGC1068            |2| 8.37e+03| 1.92e+01| 8.37e+02|Jykms|   |31| 1.14e+04| 1.14e+03|22
NGC1068            |2| 1.97e+03| 8.20e+01| 3.93e+02|Jykms|   |13| 1.15e+04| 2.34e+03| 7
NGC1068            |2| 1.13e+04| 2.20e+03| 1.70e+03|Jykms|   |  |         |         |18
NGC1068            |3| 1.16e+02| 1.40e+00| 3.48e+01|Kkms |228|22| 1.12e+04| 3.35e+03|11
NGC1068            |3| 1.68e+04| 0.00e+00| 2.95e+03|Jykms|   |43| 1.69e+04| 2.96e+03|23
NGC1068            |3| 1.71e+04| 3.40e+03| 2.56e+03|Jykms|   |  |         |         |18
NGC1056            |1| 1.12e+01| 0.00e+00| 2.80e+00|Kkms |156|24| 1.05e+02| 2.61e+01| 1
NGC1056            |2| 1.42e+01| 0.00e+00| 3.55e+00|Kkms |175|12| 2.64e+02| 6.60e+01| 1
UGC02238           |1| 6.00e+00| 0.00e+00| 1.20e+00|Kkms |288|55| 1.74e+02| 3.48e+01| 2
UGC02238           |2| 1.76e+01| 6.77e-01| 2.64e+00|Kkms |330|32| 7.96e+02| 1.23e+02| 5
UGC02238           |3| 1.87e+01| 7.16e-01| 2.80e+00|Kkms |272|22| 1.01e+03| 1.56e+02| 5
UGC02369           |1| 3.70e+00| 3.70e-01| 5.55e-01|Kkms |234|55| 1.03e+02| 1.85e+01| 8
UGC02369           |1| 1.94e+02| 3.90e+01| 2.91e+01|Jykms|   |  |         |         |18
UGC02369           |2| 9.32e+00| 3.61e-01| 1.40e+00|Kkms |230|32| 4.17e+02| 6.47e+01| 5
UGC02369           |3| 2.05e+01| 0.00e+00| 4.10e+00|Kkms |302|14| 5.12e+02| 1.02e+02|21
UGC02369           |3| 1.18e+01| 1.04e+00| 1.77e+00|Kkms |169|22| 6.35e+02| 1.10e+02| 5
UGC02369           |3| 3.87e+02| 7.70e+01| 5.80e+01|Jykms|   |  |         |         |18
NGC1222            |1| 1.74e+01| 5.24e-01| 3.47e+00|Kkms |   |21| 1.19e+02| 2.41e+01|24
NGC1222            |2| 2.88e+01| 5.60e-01| 5.75e+00|Kkms |   |10| 3.15e+02| 6.33e+01|24
NGC1222            |3| 9.80e+00| 1.32e+00| 1.47e+00|Kkms |123|22| 6.23e+02| 1.26e+02| 5
UGC02608           |1| 1.53e+01| 0.00e+00| 3.83e+00|Kkms | 87|24| 1.18e+02| 2.95e+01| 1
UGC02608           |2| 1.74e+01| 0.00e+00| 4.35e+00|Kkms | 90|12| 2.05e+02| 5.13e+01| 1
NGC1266            |1| 3.50e+01| 1.07e+00| 6.99e+00|Kkms |   |21| 1.74e+02| 3.51e+01|24
NGC1266            |1| 3.51e+01| 2.11e+00| 5.27e+00|Kkms |   |21| 1.74e+02| 2.82e+01|25
NGC1266            |2| 1.04e+02| 9.26e-01| 2.09e+01|Kkms |   |10| 5.18e+02| 1.04e+02|24
NGC1266            |2| 1.08e+02| 4.12e+00| 1.62e+01|Kkms |   |12| 6.61e+02| 1.02e+02|25
NGC1266            |3| 8.95e+02| 1.95e+01| 1.34e+02|Jykms|   |  | 8.95e+02| 1.36e+02|25
IRAS 03158+4227    |1| 2.10e+00| 0.00e+00| 7.35e-01|Kkms |180|22| 1.11e+01| 3.88e+00|17
3C 84              |1| 1.04e+02| 1.00e+00| 1.56e+01|Jykms|200|55| 9.77e+01| 1.47e+01|19
3C 84              |1| 2.50e+01| 8.00e-01| 3.75e+00|Kkms |266|21| 1.35e+02| 2.07e+01|26
3C 84              |2| 1.50e+01| 7.00e-01| 2.25e+00|Kkms |208|11| 1.00e+02| 1.57e+01|26
3C 84              |2| 3.37e+00| 6.37e-01| 5.05e-01|Kkms |166|32| 1.54e+02| 3.71e+01| 5
3C 84              |3| 9.00e+00| 8.00e-01| 2.70e+00|Kkms |248|22| 4.76e+02| 1.49e+02|11
NGC1365-SW         |1| 5.41e+01| 0.00e+00| 1.08e+01|Kkms |   |55| 1.51e+03| 3.02e+02|27
NGC1365-SW         |1| 5.78e+01| 7.40e-01| 5.78e+00|Kkms |325|55| 1.61e+03| 1.63e+02| 6
NGC1365-SW         |1| 8.96e+01| 0.00e+00| 1.79e+01|Kkms |   |44| 1.84e+03| 3.68e+02|28
NGC1365-SW         |1| 2.17e+03| 1.02e+02| 4.33e+02|Jykms|   |45| 2.12e+03| 4.35e+02| 7
NGC1365-SW         |1| 1.06e+02| 0.00e+00| 1.70e+00|Kkms |   |44| 2.18e+03| 3.49e+01| 3
NGC1365-SW         |2| 2.57e+01| 0.00e+00| 5.10e+00|Kkms |   |32| 1.43e+03| 2.84e+02|27
NGC1365-SW         |2| 1.18e+02| 0.00e+00| 2.35e+01|Kkms |   |25| 5.13e+03| 1.03e+03|28
NGC1365-SW         |3| 2.76e+02| 0.00e+00| 2.76e+01|Kkms |250|15| 2.06e+04| 2.06e+03|29
NGC1365-NE         |1| 5.78e+01| 7.40e-01| 5.78e+00|Kkms |325|55| 1.68e+03| 1.69e+02| 6
NGC1365-NE         |1| 6.22e+01| 0.00e+00| 1.24e+01|Kkms |   |55| 1.81e+03| 3.60e+02|27
NGC1365-NE         |1| 2.17e+03| 1.02e+02| 4.33e+02|Jykms|   |45| 2.13e+03| 4.38e+02| 7
NGC1365-NE         |1| 1.06e+02| 0.00e+00| 1.70e+00|Kkms |   |44| 2.18e+03| 3.50e+01| 3
NGC1365-NE         |1| 1.12e+02| 0.00e+00| 2.24e+01|Kkms |   |44| 2.31e+03| 4.61e+02|28
NGC1365-NE         |2| 3.57e+01| 0.00e+00| 7.14e+00|Kkms |   |32| 1.83e+03| 3.66e+02|27
NGC1365-NE         |2| 1.81e+02| 0.00e+00| 3.62e+01|Kkms |   |25| 6.61e+03| 1.32e+03|28
NGC1365-NE         |3| 2.77e+02| 0.00e+00| 2.76e+01|Kkms |250|15| 1.21e+04| 1.20e+03|29
NGC1482            |1| 8.10e+00| 0.00e+00| 1.62e+00|Kkms |140|55| 2.41e+02| 4.82e+01| 2
NGC1482            |1| 3.21e+01| 0.00e+00| 8.03e+00|Kkms |158|24| 2.53e+02| 6.31e+01| 1
NGC1482            |1| 2.32e+01| 0.00e+00| 5.80e+00|Kkms |259|45| 4.96e+02| 1.24e+02| 1
NGC1482            |1| 3.36e+01| 0.00e+00| 1.60e+00|Kkms |   |44| 6.92e+02| 3.29e+01| 3
NGC1482            |2| 3.34e+01| 0.00e+00| 8.35e+00|Kkms |185|12| 3.80e+02| 9.50e+01| 1
NGC1482            |2| 3.58e+01| 0.00e+00| 8.95e+00|Kkms |183|24| 1.13e+03| 2.82e+02| 1
IRAS 03521+0028    |1| 2.20e+00| 0.00e+00| 7.70e-01|Kkms |150|22| 8.73e+00| 3.06e+00|17
UGC02982           |1| 9.90e+00| 0.00e+00| 2.48e+00|Kkms |185|45| 2.04e+02| 5.10e+01| 1
UGC02982           |1| 3.56e+01| 0.00e+00| 8.90e+00|Kkms |148|24| 2.89e+02| 7.23e+01| 1
UGC02982           |2| 3.80e+01| 0.00e+00| 9.50e+00|Kkms |140|12| 5.09e+02| 1.27e+02| 1
UGC02982           |2| 1.83e+01| 0.00e+00| 4.58e+00|Kkms |178|24| 5.95e+02| 1.49e+02| 1
UGC02982           |3| 2.18e+01| 7.80e-01| 3.27e+00|Kkms |273|22| 1.42e+03| 2.18e+02| 5
IRAS04271+3849     |1| 3.41e+00| 3.86e-01| 5.11e-01|Kkms |243|55| 1.00e+02| 1.89e+01| 8
IRAS04271+3849     |2| 1.31e+01| 5.63e-01| 1.97e+00|Kkms |301|32| 5.94e+02| 9.26e+01| 5
IRAS04271+3849     |3| 1.20e+01| 6.49e-01| 1.79e+00|Kkms |251|22| 6.48e+02| 1.03e+02| 5
NGC1614            |1| 1.49e+01| 0.00e+00| 3.73e+00|Kkms | 41|24| 1.06e+02| 2.65e+01| 1
NGC1614            |1| 1.20e+01| 2.86e-01| 1.20e+00|Kkms |   |34| 1.54e+02| 1.58e+01|20
NGC1614            |1| 9.20e+00| 0.00e+00| 2.30e+00|Kkms |139|45| 1.92e+02| 4.79e+01| 1
NGC1614            |1| 3.26e+01| 5.64e-01| 6.52e+00|Kkms |   |22| 2.01e+02| 4.04e+01| 4
NGC1614            |1| 8.60e+00| 0.00e+00| 1.72e+00|Kkms |237|55| 2.53e+02| 5.07e+01| 2
NGC1614            |1| 1.52e+01| 0.00e+00| 1.10e+00|Kkms |   |44| 3.05e+02| 2.20e+01| 3
NGC1614            |1| 2.43e+02| 1.35e+01| 4.86e+01|Jykms|   |  |         |         | 7
NGC1614            |2| 3.30e+00| 0.00e+00| 8.25e-01|Kkms | 41|12| 3.06e+01| 7.66e+00| 1
NGC1614            |2| 2.99e+01| 0.00e+00| 7.47e+00|Kkms |117|24| 8.51e+02| 2.13e+02| 1
NGC1614            |2| 5.60e+01| 2.00e+00| 5.60e+00|Kkms |   |24| 1.59e+03| 1.69e+02|20
NGC1614            |3| 7.11e+01| 5.90e+00| 2.13e+01|Kkms |221|22| 3.95e+03| 1.23e+03|11
UGC03094           |1| 7.70e+00| 0.00e+00| 1.93e+00|Kkms |482|45| 1.56e+02| 3.89e+01| 1
UGC03094           |2| 1.24e+01| 0.00e+00| 3.10e+00|Kkms |113|24| 3.85e+02| 9.63e+01| 1
IRAS F05189-2524   |1| 0.00e+00| 5.10e-01| 0.00e+00|Kkms |   |55| 0.00e+00| 1.43e+01| 6
IRAS F05189-2524   |1| 2.60e+00| 0.00e+00| 5.20e-01|Kkms |   |44| 4.83e+01| 9.65e+00|12
IRAS F05189-2524   |1| 2.60e+00| 0.00e+00| 5.20e-01|Kkms |203|55| 7.28e+01| 1.46e+01| 2
IRAS F05189-2524   |1| 9.24e+01| 0.00e+00| 1.85e+01|Jykms|   |21| 1.03e+02| 2.06e+01| 7
IRAS F05189-2524   |1| 4.80e+01| 7.00e+00| 7.20e+00|Jykms|   |  |         |         |18
IRAS F05189-2524   |2| 1.30e+02| 2.20e+01| 1.95e+01|Jykms|   |  |         |         |18
IRAS F05189-2524   |3| 2.56e+02| 3.60e+01| 3.84e+01|Jykms|   |  |         |         |18
IRAS F05189-2524   |4| 0.00e+00| 6.89e+02| 0.00e+00|Jykms|   |11| 0.00e+00| 8.61e+02|18
IRAS F05189-2524   |6| 6.38e+02| 2.20e+02| 1.60e+02|Jykms|   | 8| 8.38e+02| 3.57e+02|18
SPT-S 053817-5030.8|1| 1.20e+00| 2.00e-01| 1.80e-01|Jykms|500|17| 1.36e+00| 3.05e-01|30
MCG+08-11-002      |1| 9.67e+00| 5.25e-01| 1.45e+00|Kkms |370|55| 2.88e+02| 4.60e+01| 8
MCG+08-11-002      |2| 3.00e+01| 6.26e-01| 4.50e+00|Kkms |425|32| 1.32e+03| 2.00e+02| 5
MCG+08-11-002      |3| 2.67e+01| 4.92e-01| 4.00e+00|Kkms |394|22| 1.33e+03| 2.01e+02| 5
NGC1961            |2| 3.60e+01| 4.76e-01| 5.41e+00|Kkms |401|32| 2.14e+03| 3.22e+02| 5
NGC1961            |3| 2.91e+01| 6.73e-01| 4.36e+00|Kkms |308|22| 2.83e+03| 4.29e+02| 5
UGC03351           |1| 5.58e+01| 4.80e-01| 1.12e+01|Kkms |   |22| 3.76e+02| 7.53e+01| 4
UGC03351           |1| 4.11e+02| 0.00e+00| 8.22e+01|Jykms|   |21| 5.64e+02| 1.13e+02| 7
UGC03351           |2| 5.08e+02| 3.66e+01| 1.02e+02|Jykms|   |13| 9.28e+02| 1.97e+02| 7
UGC03351           |3| 3.10e+01| 9.36e-01| 4.65e+00|Kkms |402|22| 1.88e+03| 2.88e+02| 5
IRAS05442+1732     |1| 1.46e+01| 0.00e+00| 3.65e+00|Kkms |196|24| 9.59e+01| 2.40e+01| 1
IRAS05442+1732     |1| 5.50e+00| 0.00e+00| 1.38e+00|Kkms |285|45| 1.14e+02| 2.85e+01| 1
IRAS05442+1732     |2| 2.62e+01| 0.00e+00| 6.55e+00|Kkms |220|12| 1.93e+02| 4.83e+01| 1
IRAS05442+1732     |2| 8.50e+00| 0.00e+00| 2.12e+00|Kkms |397|24| 2.23e+02| 5.58e+01| 1
IRAS05442+1732     |3| 1.63e+01| 9.25e-01| 2.44e+00|Kkms |211|22| 8.21e+02| 1.32e+02| 5
IRAS 06035-7102    |1| 1.30e+00| 0.00e+00| 2.60e-01|Kkms |   |44| 2.18e+01| 4.35e+00|12
IRAS 06035-7102    |1| 3.18e+01| 0.00e+00| 6.36e+00|Jykms|   |45| 3.18e+01| 6.36e+00| 7
NGC2146-NW         |1| 4.80e+01| 8.57e-01| 4.80e+00|Kkms |   |34| 7.20e+02| 7.31e+01|20
NGC2146-NW         |1| 8.86e+01| 0.00e+00| 2.80e+00|Kkms |   |33| 1.28e+03| 4.05e+01| 3
NGC2146-NW         |1| 1.15e+03| 2.67e+01| 2.29e+02|Jykms|   |  |         |         | 7
NGC2146-NW         |2| 1.26e+03| 1.73e+01| 2.52e+02|Jykms|   |12| 4.74e+03| 9.51e+02| 7
NGC2146-NW         |2| 1.19e+02| 1.25e+00| 1.19e+01|Kkms |   |28| 5.73e+03| 5.76e+02|20
NGC2146-NW         |3| 6.69e+01| 1.50e+00| 2.01e+01|Kkms |124|22| 5.64e+03| 1.70e+03|11
NGC2146-nuc        |1| 4.80e+01| 8.57e-01| 4.80e+00|Kkms |   |34| 6.97e+02| 7.08e+01|20
NGC2146-nuc        |1| 8.86e+01| 0.00e+00| 2.80e+00|Kkms |   |33| 1.24e+03| 3.91e+01| 3
NGC2146-nuc        |1| 1.15e+03| 2.67e+01| 2.29e+02|Jykms|   |  |         |         | 7
NGC2146-nuc        |2| 1.26e+03| 1.73e+01| 2.52e+02|Jykms|   |12| 3.64e+03| 7.30e+02| 7
NGC2146-nuc        |2| 1.19e+02| 1.25e+00| 1.19e+01|Kkms |   |28| 5.38e+03| 5.41e+02|20
NGC2146-nuc        |3| 6.69e+01| 1.50e+00| 2.01e+01|Kkms |124|22| 5.07e+03| 1.53e+03|11
NGC2146-SE         |1| 4.80e+01| 8.57e-01| 4.80e+00|Kkms |   |34| 7.18e+02| 7.29e+01|20
NGC2146-SE         |1| 8.86e+01| 0.00e+00| 2.80e+00|Kkms |   |33| 1.28e+03| 4.04e+01| 3
NGC2146-SE         |1| 1.15e+03| 2.67e+01| 2.29e+02|Jykms|   |  |         |         | 7
NGC2146-SE         |2| 1.26e+03| 1.73e+01| 2.52e+02|Jykms|   |12| 4.75e+03| 9.52e+02| 7
NGC2146-SE         |2| 4.74e+01| 9.00e-01| 4.74e+00|Kkms |   |  |         |         |20
NGC2146-SE         |3| 6.69e+01| 1.50e+00| 2.01e+01|Kkms |124|22| 5.60e+03| 1.69e+03|11
IRAS 06206-6315    |1| 2.10e+00| 0.00e+00| 4.20e-01|Kkms |   |44| 3.39e+01| 6.78e+00|12
IRAS 06206-6315    |1| 5.14e+01| 0.00e+00| 1.03e+01|Jykms|   |45| 5.12e+01| 1.02e+01| 7
ESO255-IG007       |1| 3.30e+00| 0.00e+00| 6.60e-01|Kkms |   |44| 6.15e+01| 1.23e+01|12
ESO255-IG007       |1| 7.18e+01| 1.90e+00| 1.44e+01|Jykms|   |45| 7.09e+01| 1.43e+01| 7
ESO255-IG007       |1| 3.80e+00| 1.00e-01| 3.80e-01|Kkms |182|45| 7.34e+01| 7.59e+00|13
ESO255-IG007       |2| 8.50e+00| 3.00e-01| 8.50e-01|Kkms |195|24| 2.34e+02| 2.48e+01|13
ESO255-IG007       |2| 1.74e+02| 6.20e+00| 3.48e+01|Jykms|   |  |         |         | 7
UGC03608           |2| 1.33e+01| 7.36e-01| 1.99e+00|Kkms |171|32| 6.15e+02| 9.84e+01| 5
UGC03608           |3| 1.81e+01| 1.08e+00| 2.72e+00|Kkms |199|22| 1.05e+03| 1.70e+02| 5
NGC2342a           |1| 7.10e+00| 0.00e+00| 1.77e+00|Kkms |265|45| 1.45e+02| 3.63e+01| 1
NGC2342a           |1| 2.46e+01| 0.00e+00| 6.15e+00|Kkms | 92|24| 2.53e+02| 6.32e+01| 1
NGC2342a           |2| 1.31e+01| 0.00e+00| 3.27e+00|Kkms |262|24| 5.39e+02| 1.35e+02| 1
NGC2342a           |2| 3.32e+01| 0.00e+00| 8.30e+00|Kkms |175|12| 9.30e+02| 2.32e+02| 1
NGC2369            |1| 2.37e+01| 0.00e+00| 4.74e+00|Kkms |   |44| 4.81e+02| 9.62e+01|12
NGC2369            |1| 3.71e+01| 1.43e+00| 3.71e+00|Kkms |   |34| 4.90e+02| 5.25e+01|20
NGC2369            |1| 5.54e+02| 5.70e+00| 1.11e+02|Jykms|   |45| 5.48e+02| 1.10e+02| 7
NGC2369            |1| 2.93e+01| 3.00e-01| 2.93e+00|Kkms |334|45| 6.18e+02| 6.21e+01|13
NGC2369            |1| 3.51e+01| 0.00e+00| 1.10e+00|Kkms |   |44| 7.13e+02| 2.23e+01| 3
NGC2369            |2| 4.68e+01| 7.00e-01| 4.68e+00|Kkms |339|24| 1.39e+03| 1.41e+02|13
NGC2369            |2| 3.70e+01| 1.20e+00| 3.70e+00|Kkms |   |  |         |         |20
NGC2369            |2| 9.59e+02| 1.43e+01| 1.92e+02|Jykms|   |  |         |         | 7
NGC2388a           |1| 5.11e+01| 6.24e-01| 1.02e+01|Kkms |   |22| 3.26e+02| 6.54e+01| 4
NGC2388a           |2| 2.40e+01| 3.85e-01| 3.60e+00|Kkms |270|32| 1.12e+03| 1.69e+02| 5
NGC2388a           |3| 2.19e+01| 1.03e+00| 3.28e+00|Kkms |221|22| 1.26e+03| 1.98e+02| 5
MCG+02-20-003      |1| 1.69e+01| 3.60e-01| 3.38e+00|Kkms |   |22| 1.00e+02| 2.02e+01| 4
MCG+02-20-003      |2| 5.42e+00| 5.56e-01| 8.13e-01|Kkms |234|32| 2.46e+02| 4.47e+01| 5
MCG+02-20-003      |3| 9.66e+00| 1.15e+00| 1.45e+00|Kkms |179|22| 5.17e+02| 9.90e+01| 5
IRAS 07598+6508    |1| 2.80e+00| 0.00e+00| 9.80e-01|Kkms |337|22| 1.07e+01| 3.74e+00|17
NGC2623            |1| 2.28e+01| 4.08e-01| 4.56e+00|Kkms |   |22| 1.14e+02| 2.28e+01| 4
NGC2623            |1| 4.80e+00| 0.00e+00| 9.60e-01|Kkms |255|55| 1.50e+02| 2.99e+01| 2
NGC2623            |1| 1.62e+02| 2.00e+01| 2.43e+01|Jykms|   |  | 1.62e+02| 3.15e+01|18
NGC2623            |1| 3.47e+02| 1.33e+01| 6.93e+01|Jykms|   |33| 3.47e+02| 7.06e+01| 7
NGC2623            |2| 2.67e+02| 4.00e+01| 4.00e+01|Jykms|   |  | 2.67e+02| 5.66e+01|18
NGC2623            |3| 6.14e+02| 9.20e+01| 9.21e+01|Jykms|   |  | 6.14e+02| 1.30e+02|18
IRAS 08572+3915    |1| 2.00e+00| 0.00e+00| 7.00e-01|Kkms |270|22| 9.70e+00| 3.40e+00|17
IRAS 08572+3915    |1| 1.05e+01| 1.50e+00| 1.57e+00|Jykms|   |  |         |         |18
IRAS 08572+3915    |2| 4.10e+01| 1.20e+01| 6.15e+00|Jykms|   |  |         |         |18
IRAS 08572+3915    |3| 0.00e+00| 2.40e+02| 0.00e+00|Jykms|   |  |         |         |18
IRAS 08572+3915    |6| 4.05e+02| 1.58e+02| 1.01e+02|Jykms|   | 8| 5.36e+02| 2.48e+02|18
IRAS 08572+3915    |6| 7.05e+02| 2.30e+02| 1.76e+02|Jykms|   | 8| 9.33e+02| 3.83e+02|18
NGC2764            |1| 1.62e+01| 5.80e-01| 3.24e+00|Kkms |   |21| 1.19e+02| 2.41e+01|24
NGC2764            |2| 2.44e+01| 8.47e-01| 4.88e+00|Kkms |   |10| 3.11e+02| 6.30e+01|24
NGC2798            |1| 8.10e+00| 0.00e+00| 1.90e+00|Kkms |   |33| 1.01e+02| 2.38e+01| 3
UGC05101           |1| 7.00e+01| 1.40e+01| 1.05e+01|Jykms|   |  | 7.00e+01| 1.75e+01|18
UGC05101           |1| 1.56e+01| 0.00e+00| 3.12e+00|Kkms |350|22| 7.32e+01| 1.46e+01|17
UGC05101           |1| 7.33e+01| 0.00e+00| 1.47e+01|Jykms|   |21| 7.33e+01| 1.47e+01| 7
UGC05101           |2| 3.45e+02| 6.20e+01| 5.18e+01|Jykms|   |  | 3.45e+02| 8.08e+01|18
UGC05101           |3| 5.89e+02| 9.50e+01| 8.83e+01|Jykms|   |  | 5.89e+02| 1.30e+02|18
UGC05101           |6| 0.00e+00| 4.22e+02| 0.00e+00|Jykms|   | 8| 0.00e+00| 4.22e+02|18
M82                |1| 6.67e+03| 3.35e+01| 6.67e+02|Jykms|150|45| 6.52e+03| 6.53e+02|15
M82                |1| 6.76e+02| 0.00e+00| 6.76e+01|Kkms |170|24| 7.02e+03| 7.02e+02|31
M82                |1| 4.58e+03| 0.00e+00| 9.16e+02|Jykms|   |  |         |         | 7
M82                |2| 2.86e+02| 2.20e+00| 2.86e+01|Kkms |   |30| 1.51e+04| 1.52e+03|10
M82                |2| 8.82e+02| 0.00e+00| 8.82e+01|Kkms |170|24| 3.66e+04| 3.66e+03|31
M82                |3| 5.88e+02| 0.00e+00| 5.88e+01|Kkms |170|24| 5.49e+04| 5.49e+03|31
M82                |3| 1.06e+03| 6.30e+00| 3.17e+02|Kkms |203|22| 8.93e+04| 2.68e+04|11
M82                |4| 4.46e+02| 0.00e+00| 4.46e+01|Kkms |170|24| 7.42e+04| 7.42e+03|31
M82                |6| 2.63e+02| 2.10e+01| 2.63e+01|Kkms |   |10| 5.92e+04| 7.58e+03|10
M82                |6| 2.37e+02| 0.00e+00| 2.37e+01|Kkms |170|24| 8.86e+04| 8.86e+03|31
M82                |7| 1.62e+02| 0.00e+00| 1.62e+01|Kkms |170|24| 8.26e+04| 8.26e+03|31
NGC3077            |3| 8.00e+00| 3.00e-01| 2.40e+00|Kkms | 42|22| 7.16e+02| 2.17e+02|11
NGC3110a           |1| 5.06e+01| 1.07e+01| 5.06e+00|Kkms |   |14| 2.18e+02| 5.10e+01|32
NGC3110a           |1| 3.76e+01| 5.52e-01| 7.53e+00|Kkms |   |22| 2.77e+02| 5.56e+01| 4
NGC3110a           |1| 1.30e+01| 0.00e+00| 2.60e+00|Kkms |255|55| 3.67e+02| 7.34e+01| 2
NGC3110a           |3| 3.96e+01| 8.20e+00| 3.96e+00|Kkms |   |14| 1.51e+03| 3.47e+02|32
NGC3110a           |3| 2.45e+01| 8.00e-01| 7.35e+00|Kkms |325|22| 1.62e+03| 4.90e+02|11
NGC3221            |1| 7.90e+00| 0.00e+00| 1.58e+00|Kkms |155|55| 2.09e+02| 4.18e+01| 2
NGC3221            |1| 3.35e+01| 7.10e+00| 3.35e+00|Kkms |   |14| 2.57e+02| 6.03e+01|32
NGC3221            |3| 1.69e+01| 3.50e+00| 1.69e+00|Kkms |   |14| 1.16e+03| 2.68e+02|32
NGC3227            |1| 1.47e+01| 5.30e-01| 1.47e+00|Kkms |275|55| 3.96e+02| 4.21e+01| 6
NGC3227            |3| 1.81e+01| 1.00e+00| 5.43e+00|Kkms |244|22| 1.37e+03| 4.19e+02|11
NGC3256            |1| 5.02e+01| 0.00e+00| 1.00e+01|Kkms |   |44| 1.02e+03| 2.05e+02|12
NGC3256            |1| 8.14e+01| 5.71e+00| 8.14e+00|Kkms |   |34| 1.10e+03| 1.35e+02|20
NGC3256            |1| 1.22e+03| 7.60e+00| 2.45e+02|Jykms|   |45| 1.21e+03| 2.42e+02| 7
NGC3256            |2| 3.14e+02| 8.00e+00| 3.14e+01|Kkms |   |24| 1.01e+04| 1.04e+03|20
NGC3256            |2| 2.98e+03| 1.43e+01| 5.96e+02|Jykms|   |  |         |         | 7
NGC3351            |1| 2.50e+01| 0.00e+00| 3.10e+00|Kkms |   |33| 3.33e+02| 4.13e+01| 3
NGC3351            |3| 2.60e+01| 1.40e+00| 7.80e+00|Kkms |200|22| 1.70e+03| 5.18e+02|11
IRASF10565+2448    |1| 2.20e+00| 0.00e+00| 4.40e-01|Kkms |203|55| 6.38e+01| 1.28e+01| 2
IRASF10565+2448    |1| 1.57e+01| 0.00e+00| 3.14e+00|Kkms |300|22| 7.28e+01| 1.46e+01|17
IRASF10565+2448    |1| 7.70e+01| 8.00e+00| 1.15e+01|Jykms|   |  | 7.70e+01| 1.40e+01|18
IRASF10565+2448    |1| 7.75e+01| 0.00e+00| 1.55e+01|Jykms|   |21| 7.75e+01| 1.55e+01| 7
IRASF10565+2448    |1| 3.81e+01| 8.00e+00| 3.81e+00|Kkms |   |14| 7.78e+01| 1.81e+01|32
IRASF10565+2448    |2| 3.27e+02| 3.50e+01| 4.90e+01|Jykms|   |  | 3.27e+02| 6.03e+01|18
IRASF10565+2448    |3| 2.43e+01| 5.30e+00| 2.43e+00|Kkms |   |14| 4.35e+02| 1.04e+02|32
IRASF10565+2448    |3| 2.84e+01| 0.00e+00| 5.68e+00|Kkms |187|14| 4.80e+02| 9.60e+01|21
IRASF10565+2448    |3| 1.29e+01| 2.10e+00| 1.29e+00|Kkms |   |21| 5.34e+02| 1.02e+02|10
IRASF10565+2448    |3| 5.60e+02| 5.60e+01| 8.40e+01|Jykms|   |  | 5.60e+02| 1.01e+02|18
IRASF10565+2448    |6| 5.06e+02| 1.48e+02| 1.26e+02|Jykms|   | 8| 5.06e+02| 1.95e+02|18
NGC3521            |1| 2.68e+01| 0.00e+00| 4.80e+00|Kkms |   |33| 5.25e+02| 9.41e+01| 3
NGC3521            |3| 1.45e+01| 1.40e+00| 4.35e+00|Kkms |178|22| 2.64e+03| 8.32e+02|11
NGC3627            |1| 4.48e+03| 0.00e+00| 8.95e+02|Jykms|   |  |         |         | 7
NGC3627            |2| 3.60e+03| 7.48e+01| 7.19e+02|Jykms|   |  |         |         | 7
NGC3627            |3| 2.19e+01| 9.00e-01| 6.57e+00|Kkms |142|22| 2.17e+03| 6.56e+02|11
NGC3665            |1| 1.22e+01| 6.56e-01| 2.43e+00|Kkms |   |21| 7.10e+01| 1.47e+01|24
NGC3665            |2| 1.42e+01| 8.36e-01| 2.85e+00|Kkms |   |10| 1.04e+02| 2.16e+01|24
Arp299-B           |1| 1.53e+01| 7.14e-01| 1.53e+00|Kkms |   |34| 2.45e+02| 2.71e+01|20
Arp299-B           |1| 2.93e+02| 2.67e+01| 5.87e+01|Jykms|   |33| 4.00e+02| 8.80e+01| 7
Arp299-B           |1| 5.86e+02| 1.15e+02| 8.79e+01|Jykms|   |  |         |         |18
Arp299-B           |2| 1.64e+03| 0.00e+00| 2.46e+02|Jykms|185|43| 1.64e+03| 2.46e+02|33
Arp299-B           |2| 3.12e+01| 2.08e+00| 3.12e+00|Kkms |   |28| 1.73e+03| 2.08e+02|20
Arp299-B           |3| 3.64e+01| 2.40e+00| 1.09e+01|Kkms |125|22| 3.84e+03| 1.18e+03|11
Arp299-B           |3| 8.43e+01| 0.00e+00| 1.69e+01|Kkms |167|14| 6.47e+03| 1.29e+03|21
Arp299-B           |3| 6.75e+03| 0.00e+00| 1.01e+03|Jykms|   |43| 6.74e+03| 1.01e+03|33
Arp299-B           |3| 4.36e+03| 6.55e+02| 6.54e+02|Jykms|   |  |         |         |18
Arp299-B           |4| 6.34e+03| 1.58e+03| 1.27e+03|Jykms|   |11| 3.52e+04| 1.13e+04|18
Arp299-C           |1| 1.53e+01| 7.14e-01| 1.53e+00|Kkms |   |34| 2.38e+02| 2.63e+01|20
Arp299-C           |1| 2.93e+02| 2.67e+01| 5.87e+01|Jykms|   |33| 3.88e+02| 8.52e+01| 7
Arp299-C           |1| 5.86e+02| 1.15e+02| 8.79e+01|Jykms|   |  |         |         |18
Arp299-C           |2| 2.29e+01| 2.08e+00| 2.29e+00|Kkms |   |28| 1.20e+03| 1.63e+02|20
Arp299-C           |2| 1.66e+03| 0.00e+00| 2.49e+02|Jykms| 80|43| 1.66e+03| 2.49e+02|33
Arp299-C           |3| 3.64e+01| 2.40e+00| 1.09e+01|Kkms |125|22| 3.52e+03| 1.08e+03|11
Arp299-C           |3| 8.43e+01| 0.00e+00| 1.69e+01|Kkms |167|14| 5.61e+03| 1.12e+03|21
Arp299-C           |3| 7.17e+03| 0.00e+00| 1.08e+03|Jykms|   |43| 7.16e+03| 1.07e+03|33
Arp299-C           |3| 4.36e+03| 6.55e+02| 6.54e+02|Jykms|   |  |         |         |18
Arp299-C           |4| 6.34e+03| 1.58e+03| 1.27e+03|Jykms|   |11| 2.98e+04| 9.55e+03|18
Arp299-A           |1| 1.53e+01| 7.14e-01| 1.53e+00|Kkms |   |34| 2.13e+02| 2.35e+01|20
Arp299-A           |1| 2.84e+02| 0.00e+00| 5.67e+01|Jykms|   |21| 4.43e+02| 8.85e+01| 7
Arp299-A           |1| 2.73e+01| 0.00e+00| 5.46e+00|Kkms |   |55| 7.81e+02| 1.56e+02| 2
Arp299-A           |1| 5.86e+02| 1.15e+02| 8.79e+01|Jykms|   |  |         |         |18
Arp299-A           |2| 5.38e+02| 5.40e+00| 1.08e+02|Jykms|   |13| 1.19e+03| 2.39e+02| 7
Arp299-A           |2| 1.94e+03| 0.00e+00| 2.91e+02|Jykms|325|43| 1.94e+03| 2.91e+02|33
Arp299-A           |2| 4.71e+01| 1.04e+00| 4.71e+00|Kkms |   |28| 2.00e+03| 2.05e+02|20
Arp299-A           |3| 7.91e+01| 0.00e+00| 1.58e+01|Kkms |261|14| 3.08e+03| 6.17e+02|21
Arp299-A           |3| 4.87e+01| 1.90e+00| 1.46e+01|Kkms |239|22| 3.38e+03| 1.02e+03|11
Arp299-A           |3| 8.44e+03| 0.00e+00| 1.27e+03|Jykms|   |43| 8.44e+03| 1.27e+03|33
Arp299-A           |3| 4.36e+03| 6.55e+02| 6.54e+02|Jykms|   |  |         |         |18
Arp299-A           |4| 6.34e+03| 1.58e+03| 1.27e+03|Jykms|   |11| 1.59e+04| 5.10e+03|18
ESO 320-G030       |1| 9.20e+00| 0.00e+00| 1.84e+00|Kkms |   |44| 1.87e+02| 3.74e+01|12
ESO 320-G030       |1| 2.25e+02| 0.00e+00| 4.51e+01|Jykms|   |45| 2.24e+02| 4.48e+01| 7
NGC3982            |1| 5.48e+00| 3.70e-01| 5.48e-01|Kkms |137|55| 1.49e+02| 1.80e+01|34
NGC3982            |3| 6.70e+00| 7.00e-01| 2.01e+00|Kkms | 61|22| 7.14e+02| 2.27e+02|11
NGC4038            |1| 2.31e+01| 0.00e+00| 4.63e+00|Kkms |   |43| 4.65e+02| 9.30e+01|35
NGC4038            |1| 3.00e+01| 2.86e+00| 3.00e+00|Kkms |   |34| 5.05e+02| 6.97e+01|20
NGC4038            |1| 6.76e+02| 3.39e+01| 6.76e+01|Jykms|180|45| 6.47e+02| 7.24e+01|15
NGC4038            |2| 5.10e+01| 1.00e+00| 5.10e+00|Kkms |   |  |         |         |20
NGC4038            |3| 1.50e+01| 3.20e-01| 2.26e+00|Kkms |   |43| 2.72e+03| 4.13e+02|35
NGC4038            |3| 4.40e+01| 1.00e+00| 1.32e+01|Kkms | 87|22| 4.38e+03| 1.32e+03|11
NGC4038overlap     |1| 4.39e+01| 5.71e-01| 4.39e+00|Kkms |   |34| 6.92e+02| 6.98e+01|20
NGC4038overlap     |1| 4.23e+01| 0.00e+00| 8.47e+00|Kkms |   |43| 8.47e+02| 1.69e+02|35
NGC4038overlap     |2| 5.10e+01| 1.00e+00| 5.10e+00|Kkms |   |  |         |         |20
NGC4038overlap     |3| 2.87e+01| 4.10e-01| 4.31e+00|Kkms |   |43| 5.18e+03| 7.80e+02|35
NGC4038overlap     |3| 8.26e+01| 2.30e+00| 2.48e+01|Kkms |166|22| 8.02e+03| 2.42e+03|11
NGC4051            |1| 8.82e+00| 2.80e-01| 8.82e-01|Kkms |140|55| 2.08e+02| 2.18e+01| 6
NGC4051            |2| 1.80e+01| 5.93e-01| 2.70e+00|Kkms |142|32| 1.12e+03| 1.72e+02| 5
NGC4051            |3| 1.24e+01| 7.56e-01| 1.86e+00|Kkms |142|22| 1.13e+03| 1.83e+02| 5
NGC4194            |1| 4.10e+00| 0.00e+00| 8.20e-01|Kkms |183|55| 1.22e+02| 2.45e+01| 2
NGC4194            |1| 1.65e+01| 0.00e+00| 4.12e+00|Kkms |149|24| 1.24e+02| 3.10e+01| 1
NGC4194            |1| 1.20e+01| 0.00e+00| 1.80e+00|Kkms |   |33| 1.51e+02| 2.27e+01| 3
NGC4194            |2| 5.27e+01| 0.00e+00| 1.32e+01|Kkms |170|12| 5.38e+02| 1.35e+02| 1
NGC4194            |3| 4.82e+00| 9.06e-01| 7.23e-01|Kkms |157|22| 2.84e+02| 6.82e+01| 5
NGC4254            |3| 2.40e+01| 1.70e+00| 7.20e+00|Kkms |140|22| 2.93e+03| 9.04e+02|11
NGC4321            |3| 5.69e+01| 4.20e+00| 1.71e+01|Kkms |177|22| 4.57e+03| 1.41e+03|11
NGC4388            |1| 7.92e+00| 3.70e-01| 7.92e-01|Kkms |250|55| 2.10e+02| 2.31e+01| 6
NGC4388            |2| 1.88e+01| 5.28e-01| 2.82e+00|Kkms |256|32| 1.08e+03| 1.65e+02| 5
NGC4388            |3| 1.29e+01| 7.58e-01| 1.94e+00|Kkms |238|22| 1.13e+03| 1.82e+02| 5
NGC4536            |1| 2.02e+01| 0.00e+00| 2.60e+00|Kkms |   |33| 2.73e+02| 3.51e+01| 3
TOL1238-364        |1| 2.60e+00| 0.00e+00| 6.50e-01|Kkms | 82|45| 5.43e+01| 1.36e+01| 1
TOL1238-364        |2| 8.90e+00| 0.00e+00| 2.23e+00|Kkms |170|24| 3.58e+02| 8.95e+01| 1
NGC4631            |1| 1.17e+03| 0.00e+00| 2.33e+02|Jykms|   |  |         |         | 7
NGC4631            |3| 1.77e+01| 7.00e-01| 5.31e+00|Kkms | 71|22| 2.26e+03| 6.83e+02|11
NGC4710            |1| 3.17e+01| 9.23e-01| 6.34e+00|Kkms |   |21| 2.23e+02| 4.50e+01|24
NGC4710            |2| 4.01e+01| 7.66e-01| 8.03e+00|Kkms |   |10| 4.29e+02| 8.62e+01|24
NGC4710            |3| 1.87e+01| 2.50e+00| 5.61e+00|Kkms |158|22| 1.21e+03| 3.99e+02|11
NGC4736            |3| 2.13e+01| 2.00e+00| 6.39e+00|Kkms |122|22| 2.71e+03| 8.51e+02|11
NGC4736            |3| 3.20e+01| 2.30e+00| 3.20e+00|Kkms |   |21| 4.05e+03| 4.99e+02|10
Mrk 231            |1| 1.60e+00| 0.00e+00| 3.20e-01|Kkms |167|55| 4.66e+01| 9.31e+00| 2
Mrk 231            |1| 8.80e+01| 9.00e+00| 1.32e+01|Jykms|   |  | 8.80e+01| 1.60e+01|18
Mrk 231            |1| 8.99e+01| 1.01e+01| 8.19e+00|Jykms|200|45| 8.99e+01| 1.30e+01|15
Mrk 231            |1| 1.74e+01| 0.00e+00| 4.35e+00|Kkms |186|24| 9.64e+01| 2.41e+01| 1
Mrk 231            |1| 3.40e+00| 3.20e-01| 3.40e-01|Kkms |230|55| 9.91e+01| 1.36e+01| 6
Mrk 231            |1| 2.20e+01| 0.00e+00| 4.40e+00|Kkms |230|22| 1.02e+02| 2.05e+01|17
Mrk 231            |1| 1.04e+02| 0.00e+00| 2.07e+01|Jykms|   |  | 1.04e+02| 2.07e+01| 7
Mrk 231            |2| 5.16e+01| 0.00e+00| 1.29e+01|Kkms |194|12| 2.86e+02| 7.15e+01| 1
Mrk 231            |2| 3.15e+02| 3.00e+01| 4.72e+01|Jykms|   |  | 3.15e+02| 5.60e+01|18
Mrk 231            |2| 1.19e+01| 5.00e-01| 1.19e+00|Kkms |   |30| 4.26e+02| 4.62e+01|10
Mrk 231            |3| 8.70e+00| 7.00e-01| 8.70e-01|Kkms |   |21| 3.61e+02| 4.64e+01|10
Mrk 231            |3| 5.68e+02| 8.00e+01| 8.52e+01|Jykms|   |  | 5.68e+02| 1.17e+02|18
Mrk 231            |4| 1.13e+03| 2.65e+02| 2.25e+02|Jykms|   |11| 1.13e+03| 3.48e+02|18
Mrk 231            |6| 1.32e+03| 4.00e+02| 3.30e+02|Jykms|   | 8| 1.32e+03| 5.19e+02|18
NGC4826            |1| 4.90e+01| 2.33e+00| 4.90e+00|Kkms |   |33| 7.36e+02| 8.15e+01|20
NGC4826            |1| 2.17e+03| 0.00e+00| 4.35e+02|Jykms|   |22| 4.30e+03| 8.59e+02| 7
NGC4826            |2| 5.21e+01| 2.08e+00| 5.21e+00|Kkms |   |28| 2.66e+03| 2.86e+02|20
NGC4826            |3| 8.68e+01| 5.20e+00| 2.60e+01|Kkms |214|22| 8.10e+03| 2.48e+03|11
ESO507-G070        |1| 5.80e+00| 0.00e+00| 1.16e+00|Kkms |   |44| 1.15e+02| 2.29e+01|12
ESO507-G070        |1| 1.42e+02| 0.00e+00| 2.84e+01|Jykms|   |45| 1.41e+02| 2.83e+01| 7
ESO507-G070        |1| 1.52e+02| 3.00e+01| 2.28e+01|Jykms|   |  |         |         |18
ESO507-G070        |3| 4.38e+01| 0.00e+00| 8.76e+00|Kkms |479|14| 9.51e+02| 1.90e+02|21
ESO507-G070        |3| 8.64e+02| 1.73e+02| 1.30e+02|Jykms|   |  |         |         |18
NGC5055            |1| 4.11e+01| 0.00e+00| 1.50e+00|Kkms |   |33| 6.91e+02| 2.52e+01| 3
NGC5055            |1| 4.33e+01| 3.33e+00| 4.33e+00|Kkms |   |33| 7.29e+02| 9.19e+01|20
NGC5055            |1| 4.69e+03| 0.00e+00| 9.38e+02|Jykms|   |22| 1.14e+04| 2.28e+03| 7
NGC5055            |3| 2.58e+01| 3.50e+00| 7.74e+00|Kkms |190|22| 2.95e+03| 9.71e+02|11
Arp193             |1| 0.00e+00| 4.90e+00| 0.00e+00|Jykms|   |55| 0.00e+00| 4.67e+00|19
Arp193             |1| 4.10e+00| 0.00e+00| 1.20e+00|Kkms |   |33| 4.77e+01| 1.40e+01| 3
Arp193             |1| 2.40e+00| 0.00e+00| 4.80e-01|Kkms |267|55| 7.02e+01| 1.40e+01| 2
Arp193             |1| 1.71e+02| 0.00e+00| 3.42e+01|Jykms|   |21| 2.00e+02| 3.99e+01| 7
Arp193             |1| 3.60e+01| 0.00e+00| 7.20e+00|Kkms |410|22| 2.04e+02| 4.08e+01|17
Arp193             |1| 9.06e+01| 1.84e+01| 9.06e+00|Kkms |   |14| 2.52e+02| 5.70e+01|32
Arp193             |1| 1.94e+02| 1.60e+01| 2.91e+01|Jykms|   |  |         |         |18
Arp193             |2| 1.30e+01| 5.77e-01| 1.95e+00|Kkms |290|32| 5.72e+02| 8.95e+01| 5
Arp193             |2| 8.50e+02| 1.30e+02| 1.28e+02|Jykms|   |  |         |         |18
Arp193             |3| 2.05e+01| 1.70e+00| 6.15e+00|Kkms |240|22| 1.05e+03| 3.25e+02|11
Arp193             |3| 6.33e+01| 1.29e+01| 6.33e+00|Kkms |   |14| 1.55e+03| 3.51e+02|32
Arp193             |3| 1.29e+03| 1.71e+02| 1.94e+02|Jykms|   |  |         |         |18
Arp193             |6| 0.00e+00| 6.30e+02| 0.00e+00|Jykms|   | 8| 0.00e+00| 9.41e+02|18
NGC5104            |1| 6.20e+00| 0.00e+00| 1.55e+00|Kkms |361|45| 1.28e+02| 3.21e+01| 1
NGC5104            |1| 6.26e+01| 1.27e+01| 6.26e+00|Kkms |   |14| 1.70e+02| 3.84e+01|32
NGC5104            |1| 1.50e+02| 3.00e+01| 2.25e+01|Jykms|   |  |         |         |18
NGC5104            |2| 1.30e+01| 6.91e-01| 1.94e+00|Kkms |405|32| 5.79e+02| 9.23e+01| 5
NGC5104            |3| 1.28e+01| 7.95e-01| 1.92e+00|Kkms |276|22| 6.55e+02| 1.06e+02| 5
NGC5104            |3| 3.36e+01| 6.80e+00| 3.36e+00|Kkms |   |14| 7.99e+02| 1.80e+02|32
NGC5104            |3| 7.06e+02| 1.43e+02| 1.06e+02|Jykms|   |  |         |         |18
Cen A              |1| 6.90e+01| 0.00e+00| 1.38e+01|Kkms |   |44| 1.43e+03| 2.85e+02|36
Cen A              |1| 7.10e+01| 4.00e+00| 7.10e+00|Kkms |   |45| 1.50e+03| 1.72e+02|37
Cen A              |2| 7.00e+01| 7.00e+00| 7.00e+00|Kkms |   |22| 2.97e+03| 4.20e+02|37
Cen A              |3| 1.30e+02| 0.00e+00| 2.99e+01|Kkms |150|21| 1.18e+04| 2.72e+03|38
NGC5135            |1| 1.11e+01| 0.00e+00| 2.22e+00|Kkms | 76|55| 3.25e+02| 6.49e+01| 2
NGC5135            |1| 1.50e+01| 7.00e-01| 1.50e+00|Kkms |100|55| 4.39e+02| 4.85e+01| 6
NGC5135            |1| 4.26e+02| 0.00e+00| 8.53e+01|Jykms|   |22| 5.26e+02| 1.05e+02| 7
NGC5135            |1| 3.82e+02| 4.80e+01| 5.73e+01|Jykms|   |  |         |         |18
NGC5135            |2| 1.24e+03| 1.20e+02| 1.85e+02|Jykms|   |  |         |         |18
NGC5135            |3| 1.96e+03| 2.95e+02| 2.94e+02|Jykms|   |  |         |         |18
NGC5194            |1| 3.74e+01| 4.14e+00| 5.61e+00|Kkms |125|55| 8.90e+02| 1.66e+02| 8
NGC5194            |2| 4.86e+01| 6.03e-01| 7.30e+00|Kkms | 96|32| 3.56e+03| 5.36e+02| 5
NGC5194            |3| 4.44e+01| 2.80e+00| 1.33e+01|Kkms | 61|22| 7.06e+03| 2.16e+03|11
NGC5194            |4| 3.67e+01| 2.40e+00| 3.67e+00|Kkms |   |14| 1.19e+04| 1.43e+03|10
IC4280             |1| 1.15e+01| 0.00e+00| 2.88e+00|Kkms |153|45| 2.38e+02| 5.96e+01| 1
IC4280             |1| 3.23e+01| 0.00e+00| 8.07e+00|Kkms |152|24| 2.64e+02| 6.60e+01| 1
IC4280             |2| 4.66e+01| 0.00e+00| 1.17e+01|Kkms |148|12| 6.89e+02| 1.72e+02| 1
M83                |1| 2.05e+03| 0.00e+00| 2.05e+02|Jykms|100|45| 1.99e+03| 1.99e+02|15
M83                |1| 6.54e+02| 3.33e+01| 1.31e+02|Jykms|   |  |         |         | 7
M83                |3| 1.26e+02| 0.00e+00| 2.90e+01|Kkms | 94|21| 1.17e+04| 2.69e+03|38
M83                |3| 1.54e+02| 3.10e+00| 4.62e+01|Kkms |112|22| 1.47e+04| 4.42e+03|11
Mrk 273            |1| 4.33e+01| 1.49e+01| 4.33e+00|Jykms|   |45| 4.30e+01| 1.55e+01|15
Mrk 273            |1| 2.30e+00| 0.00e+00| 4.60e-01|Kkms |122|55| 6.44e+01| 1.29e+01| 2
Mrk 273            |1| 1.90e+01| 0.00e+00| 3.80e+00|Kkms |300|22| 1.03e+02| 2.06e+01|17
Mrk 273            |1| 1.98e+01| 0.00e+00| 4.95e+00|Kkms |244|24| 1.25e+02| 3.13e+01| 1
Mrk 273            |1| 9.73e+01| 0.00e+00| 1.95e+01|Jykms|   |  |         |         | 7
Mrk 273            |1| 8.20e+01| 9.00e+00| 1.23e+01|Jykms|   |  |         |         |18
Mrk 273            |2| 1.98e+01| 0.00e+00| 4.95e+00|Kkms |201|12| 1.52e+02| 3.81e+01| 1
Mrk 273            |2| 2.70e+02| 3.50e+01| 4.05e+01|Jykms|   |  |         |         |18
Mrk 273            |3| 4.82e+02| 8.20e+01| 7.23e+01|Jykms|   |  |         |         |18
Mrk 273            |6| 4.88e+02| 1.56e+02| 1.22e+02|Jykms|   | 8| 7.50e+02| 3.04e+02|18
4C 12.50           |1| 8.00e+00| 4.00e-01| 1.20e+00|Jykms|400|55| 7.48e+00| 1.18e+00|19
UGC08739           |1| 4.42e+01| 9.00e+00| 4.42e+00|Kkms |   |14| 2.61e+02| 5.91e+01|32
UGC08739           |1| 1.18e+02| 2.40e+01| 1.77e+01|Jykms|   |  |         |         |18
UGC08739           |2| 2.62e+00| 2.42e-01| 3.93e-01|Kkms |258|32| 1.32e+02| 2.32e+01| 5
UGC08739           |3| 4.83e+01| 9.90e+00| 4.83e+00|Kkms |   |14| 2.55e+03| 5.81e+02|32
UGC08739           |3| 1.13e+03| 2.31e+02| 1.69e+02|Jykms|   |  |         |         |18
OQ 208             |1| 0.00e+00| 7.90e+00| 0.00e+00|Jykms|   |55| 0.00e+00| 7.44e+00|19
NGC5653            |1| 5.30e+00| 0.00e+00| 1.06e+00|Kkms |206|55| 1.52e+02| 3.04e+01| 2
NGC5653            |1| 9.90e+00| 0.00e+00| 2.48e+00|Kkms | 88|45| 2.07e+02| 5.19e+01| 1
NGC5653            |1| 6.11e+01| 1.26e+01| 6.11e+00|Kkms |   |14| 3.19e+02| 7.32e+01|32
NGC5653            |1| 4.39e+01| 6.84e-01| 8.77e+00|Kkms |   |22| 3.44e+02| 6.90e+01| 4
NGC5653            |1| 1.87e+02| 2.70e+01| 2.81e+01|Jykms|   |  |         |         |18
NGC5653            |3| 3.84e+01| 7.70e+00| 3.84e+00|Kkms |   |14| 1.79e+03| 4.00e+02|32
NGC5653            |3| 8.06e+02| 1.62e+02| 1.21e+02|Jykms|   |  |         |         |18
IRAS 14348-1447    |1| 1.70e+00| 0.00e+00| 3.40e-01|Kkms |   |44| 2.82e+01| 5.64e+00|12
IRAS 14348-1447    |1| 4.16e+01| 0.00e+00| 8.32e+00|Jykms|   |45| 4.14e+01| 8.28e+00| 7
IRAS 14348-1447    |1| 1.70e+00| 0.00e+00| 3.40e-01|Kkms |198|55| 4.24e+01| 8.48e+00| 2
IRAS 14348-1447    |1| 5.60e+01| 8.00e+00| 8.40e+00|Jykms|   |  |         |         |18
IRAS 14348-1447    |2| 2.12e+02| 3.50e+01| 3.18e+01|Jykms|   |  |         |         |18
IRAS 14348-1447    |3| 1.94e+01| 0.00e+00| 3.88e+00|Kkms |240|14| 3.37e+02| 6.73e+01|21
IRAS 14348-1447    |3| 3.60e+02| 6.70e+01| 5.40e+01|Jykms|   |  |         |         |18
NGC5713            |1| 1.64e+01| 4.10e+00| 1.64e+00|Kkms |   |14| 1.26e+02| 3.40e+01|32
NGC5713            |1| 2.11e+01| 0.00e+00| 5.28e+00|Kkms |104|45| 4.43e+02| 1.11e+02| 1
NGC5713            |1| 5.42e+01| 0.00e+00| 1.36e+01|Kkms |100|24| 5.98e+02| 1.49e+02| 1
NGC5713            |1| 5.06e+02| 0.00e+00| 1.01e+02|Jykms|   |22| 1.00e+03| 2.01e+02| 7
NGC5713            |2| 3.80e+01| 0.00e+00| 9.50e+00|Kkms | 95|24| 1.68e+03| 4.19e+02| 1
NGC5713            |2| 7.62e+01| 0.00e+00| 1.91e+01|Kkms |101|12| 2.15e+03| 5.37e+02| 1
NGC5713            |3| 2.72e+01| 5.50e+00| 2.72e+00|Kkms |   |14| 1.87e+03| 4.22e+02|32
IRAS 14378-3651    |1| 2.45e+01| 0.00e+00| 4.90e+00|Jykms|   |45| 2.45e+01| 4.90e+00| 7
3C 305             |1| 0.00e+00| 8.60e+00| 0.00e+00|Jykms|   |55| 0.00e+00| 8.00e+00|19
VV340a             |1| 7.12e+00| 4.00e-01| 1.07e+00|Kkms |543|55| 1.95e+02| 3.12e+01| 8
VV340a             |3| 5.20e+00| 1.70e+00| 5.20e-01|Kkms |   |14| 1.35e+02| 4.63e+01|32
VV340a             |3| 1.81e+01| 1.10e+00| 5.43e+00|Kkms |548|22| 9.57e+02| 2.93e+02|11
VV340a             |3| 4.81e+01| 0.00e+00| 9.62e+00|Kkms |502|14| 1.19e+03| 2.39e+02|21
NGC5866            |1| 6.33e+00| 4.35e-01| 9.50e-01|Kkms |369|55| 1.83e+02| 3.02e+01| 8
NGC5866            |3| 0.00e+00| 8.60e+00| 0.00e+00|Kkms |200|22| 0.00e+00| 6.63e+02|11
NGC5866            |3| 7.95e+00| 5.80e-01| 1.19e+00|Kkms |260|22| 6.13e+02| 1.02e+02| 5
CGCG049-057        |1| 2.74e+01| 6.00e+00| 2.74e+00|Kkms |   |14| 6.11e+01| 1.47e+01|32
CGCG049-057        |1| 3.40e+00| 0.00e+00| 6.80e-01|Kkms |230|55| 1.08e+02| 2.15e+01| 2
CGCG049-057        |1| 1.18e+02| 0.00e+00| 2.36e+01|Jykms|   |21| 1.18e+02| 2.36e+01| 7
CGCG049-057        |1| 1.20e+02| 1.10e+01| 1.80e+01|Jykms|   |  | 1.20e+02| 2.11e+01|18
CGCG049-057        |2| 3.56e+02| 4.60e+00| 7.13e+01|Jykms|   |13| 3.56e+02| 7.14e+01| 7
CGCG049-057        |2| 1.21e+01| 9.96e-01| 1.82e+00|Kkms |249|32| 5.19e+02| 8.87e+01| 5
CGCG049-057        |2| 6.05e+02| 9.20e+01| 9.08e+01|Jykms|   |  | 6.05e+02| 1.29e+02|18
CGCG049-057        |3| 2.28e+01| 4.90e+00| 2.28e+00|Kkms |   |14| 4.45e+02| 1.06e+02|32
CGCG049-057        |3| 7.10e+02| 1.00e+02| 1.06e+02|Jykms|   |  | 7.10e+02| 1.46e+02|18
CGCG049-057        |4| 1.12e+03| 2.62e+02| 2.24e+02|Jykms|   |11| 1.12e+03| 3.45e+02|18
CGCG049-057        |6| 9.04e+02| 2.41e+02| 2.26e+02|Jykms|   | 8| 9.04e+02| 3.30e+02|18
VV705              |1| 8.30e+00| 0.00e+00| 2.08e+00|Kkms | 93|24| 5.17e+01| 1.29e+01| 1
VV705              |1| 2.00e+00| 0.00e+00| 4.00e-01|Kkms |170|55| 5.57e+01| 1.11e+01| 2
VV705              |1| 1.14e+02| 2.30e+01| 1.71e+01|Jykms|   |  |         |         |18
VV705              |2| 1.45e+01| 0.00e+00| 3.62e+00|Kkms |110|12| 1.06e+02| 2.66e+01| 1
VV705              |3| 4.20e+00| 4.00e-01| 1.26e+00|Kkms | 88|22| 2.02e+02| 6.35e+01|11
VV705              |3| 1.46e+01| 3.30e+00| 1.46e+00|Kkms |   |14| 3.32e+02| 8.22e+01|32
VV705              |3| 1.99e+01| 0.00e+00| 3.98e+00|Kkms |121|14| 4.31e+02| 8.62e+01|21
VV705              |3| 3.64e+02| 7.30e+01| 5.46e+01|Jykms|   |  |         |         |18
IRAS 15250+3609    |3| 1.03e+01| 3.30e+00| 1.03e+00|Kkms |   |14| 1.78e+02| 5.97e+01|32
NGC5936            |1| 5.70e+00| 0.00e+00| 1.14e+00|Kkms |155|55| 1.62e+02| 3.23e+01| 2
NGC5936            |1| 3.29e+01| 3.60e-01| 6.59e+00|Kkms |   |22| 2.50e+02| 5.01e+01| 4
NGC5936            |1| 5.64e+01| 1.18e+01| 5.64e+00|Kkms |   |14| 2.57e+02| 5.96e+01|32
NGC5936            |2| 1.47e+01| 8.43e-01| 2.21e+00|Kkms |162|32| 7.44e+02| 1.19e+02| 5
NGC5936            |3| 3.78e+01| 7.60e+00| 3.78e+00|Kkms |   |14| 1.52e+03| 3.42e+02|32
NGC5936            |3| 2.60e+01| 1.26e+00| 3.90e+00|Kkms |160|22| 1.78e+03| 2.80e+02| 5
Arp220             |1| 9.40e+00| 0.00e+00| 1.88e+00|Kkms |360|55| 2.80e+02| 5.61e+01| 2
Arp220             |1| 1.26e+02| 2.62e+01| 1.26e+01|Kkms |   |14| 3.30e+02| 7.59e+01|32
Arp220             |1| 4.02e+02| 0.00e+00| 2.23e+01|Jykms|420|45| 4.00e+02| 2.21e+01|15
Arp220             |1| 1.09e+02| 0.00e+00| 2.18e+01|Kkms |480|22| 6.02e+02| 1.20e+02|17
Arp220             |1| 2.05e+01| 8.20e-01| 2.05e+00|Kkms |470|55| 6.12e+02| 6.59e+01| 6
Arp220             |1| 4.19e+02| 3.60e+01| 6.28e+01|Jykms|   |  |         |         |18
Arp220             |1| 5.15e+02| 0.00e+00| 1.03e+02|Jykms|   |  |         |         | 7
Arp220             |2| 1.55e+03| 3.11e+02| 0.00e+00|Jykms|420|20| 1.73e+03| 3.48e+02|39
Arp220             |2| 6.51e+02| 3.24e+01| 1.30e+02|Jykms|   |  |         |         | 7
Arp220             |2| 1.13e+03| 6.90e+01| 1.69e+02|Jykms|   |  |         |         |18
Arp220             |3| 2.79e+01| 1.90e+00| 2.79e+00|Kkms |   |21| 1.38e+03| 1.67e+02|10
Arp220             |3| 7.42e+01| 1.49e+01| 7.42e+00|Kkms |   |14| 1.70e+03| 3.81e+02|32
Arp220             |3| 5.85e+01| 1.90e+00| 1.76e+01|Kkms |379|22| 2.91e+03| 8.78e+02|11
Arp220             |3| 3.17e+03| 6.34e+02| 0.00e+00|Jykms|510|14| 3.79e+03| 7.59e+02|39
Arp220             |3| 3.67e+03| 4.05e+02| 5.51e+02|Jykms|   |  |         |         |18
Arp220             |6| 3.13e+03| 8.10e+02| 7.82e+02|Jykms|   | 8| 4.08e+03| 1.47e+03|18
NGC5990            |1| 1.04e+01| 0.00e+00| 2.60e+00|Kkms |350|45| 2.18e+02| 5.46e+01| 1
NGC5990            |1| 3.67e+01| 0.00e+00| 9.18e+00|Kkms |232|24| 2.80e+02| 6.99e+01| 1
NGC5990            |1| 8.67e+01| 2.00e+01| 8.67e+00|Kkms |   |14| 3.20e+02| 8.04e+01|32
NGC5990            |1| 2.24e+02| 5.20e+01| 3.36e+01|Jykms|   |  |         |         |18
NGC5990            |2| 8.20e+00| 0.00e+00| 2.05e+00|Kkms |295|24| 2.50e+02| 6.25e+01| 1
NGC5990            |2| 3.06e+01| 0.00e+00| 7.65e+00|Kkms |202|12| 3.43e+02| 8.57e+01| 1
NGC5990            |3| 2.81e+01| 5.90e+00| 2.81e+00|Kkms |   |14| 9.15e+02| 2.13e+02|32
NGC5990            |3| 3.42e+01| 2.67e+00| 5.14e+00|Kkms |304|22| 2.06e+03| 3.48e+02| 5
NGC5990            |3| 6.36e+02| 1.33e+02| 9.54e+01|Jykms|   |  |         |         |18
NGC6052            |1| 1.64e+01| 0.00e+00| 4.10e+00|Kkms |123|24| 1.36e+02| 3.39e+01| 1
NGC6052            |1| 3.06e+01| 8.00e+00| 3.06e+00|Kkms |   |14| 1.40e+02| 3.92e+01|32
NGC6052            |2| 2.47e+01| 0.00e+00| 6.17e+00|Kkms |122|12| 3.69e+02| 9.22e+01| 1
NGC6052            |3| 1.78e+01| 3.70e+00| 1.78e+00|Kkms |   |14| 7.22e+02| 1.67e+02|32
CGCG052-037        |1| 2.64e+01| 6.30e+00| 2.64e+00|Kkms |   |14| 7.31e+01| 1.89e+01|32
CGCG052-037        |1| 6.30e+01| 1.50e+01| 9.45e+00|Jykms|   |  |         |         |18
CGCG052-037        |2| 1.34e+01| 6.77e-01| 2.00e+00|Kkms |282|32| 5.86e+02| 9.28e+01| 5
CGCG052-037        |3| 2.76e+01| 5.70e+00| 2.76e+00|Kkms |   |14| 6.71e+02| 1.54e+02|32
CGCG052-037        |3| 1.85e+01| 1.70e+00| 2.77e+00|Kkms |260|22| 9.39e+02| 1.65e+02| 5
CGCG052-037        |3| 5.80e+02| 1.20e+02| 8.70e+01|Jykms|   |  |         |         |18
NGC6156            |1| 1.38e+01| 0.00e+00| 3.45e+00|Kkms |182|45| 2.86e+02| 7.15e+01| 1
NGC6156            |1| 1.60e+01| 0.00e+00| 7.00e-01|Kkms |   |44| 3.23e+02| 1.41e+01| 3
NGC6156            |2| 3.08e+01| 0.00e+00| 7.70e+00|Kkms |213|24| 1.39e+03| 3.48e+02| 1
ESO069-IG006       |1| 7.30e+00| 0.00e+00| 1.46e+00|Kkms |   |44| 1.34e+02| 2.68e+01|12
ESO069-IG006       |1| 1.79e+02| 0.00e+00| 3.58e+01|Jykms|   |45| 1.78e+02| 3.56e+01| 7
IRASF16399-0937    |1| 1.18e+02| 0.00e+00| 2.36e+01|Jykms|   |21| 1.59e+02| 3.17e+01| 7
IRASF16399-0937    |2| 6.74e+01| 9.20e+00| 1.35e+01|Jykms|   |13| 1.13e+02| 2.73e+01| 7
IRASF16399-0937    |3| 1.11e+01| 1.00e+00| 1.66e+00|Kkms |240|22| 6.37e+02| 1.12e+02| 5
NGC6240            |1| 2.39e+02| 1.64e+01| 2.39e+01|Jykms|420|45| 2.36e+02| 2.87e+01|15
NGC6240            |1| 9.00e+00| 0.00e+00| 1.80e+00|Kkms |280|55| 2.57e+02| 5.14e+01| 2
NGC6240            |1| 6.90e+01| 0.00e+00| 1.38e+01|Kkms |370|22| 4.16e+02| 8.32e+01|17
NGC6240            |1| 3.33e+02| 0.00e+00| 6.66e+01|Jykms|   |  |         |         | 7
NGC6240            |1| 3.22e+02| 2.90e+01| 4.83e+01|Jykms|   |  |         |         |18
NGC6240            |2| 1.74e+03| 3.50e+02| 0.00e+00|Jykms|410|20| 2.19e+03| 4.39e+02|39
NGC6240            |2| 4.57e+02| 1.25e+01| 9.14e+01|Jykms|   |  |         |         | 7
NGC6240            |2| 1.49e+03| 2.53e+02| 2.24e+02|Jykms|   |  |         |         |18
NGC6240            |3| 7.49e+01| 2.20e+00| 2.25e+01|Kkms |355|22| 4.06e+03| 1.22e+03|11
NGC6240            |3| 3.20e+03| 6.42e+02| 0.00e+00|Jykms|390|14| 4.65e+03| 9.32e+02|39
NGC6240            |3| 3.20e+03| 6.42e+02| 4.81e+02|Jykms|   |  |         |         |18
NGC6240            |6| 3.32e+03| 8.60e+02| 8.30e+02|Jykms|   | 8| 5.87e+03| 2.11e+03|18
IRASF16516-0948    |1| 2.96e+00| 2.26e-01| 4.44e-01|Kkms |283|55| 7.94e+01| 1.34e+01| 8
IRASF16516-0948    |2| 1.52e+01| 3.09e-01| 2.29e+00|Kkms |289|32| 7.58e+02| 1.15e+02| 5
IRASF16516-0948    |3| 1.36e+01| 1.16e+00| 2.04e+00|Kkms |211|22| 9.29e+02| 1.60e+02| 5
NGC6286a           |1| 6.80e+00| 0.00e+00| 1.36e+00|Kkms |440|55| 1.94e+02| 3.89e+01| 2
NGC6286a           |2| 1.32e+01| 4.54e-01| 1.98e+00|Kkms |319|32| 6.27e+02| 9.65e+01| 5
NGC6286a           |3| 1.33e+01| 1.80e+00| 3.99e+00|Kkms |282|22| 8.34e+02| 2.74e+02|11
IRASF17138-1017    |1| 3.28e+01| 4.20e-01| 6.57e+00|Kkms |   |22| 1.95e+02| 3.91e+01| 4
IRASF17138-1017    |2| 2.23e+01| 8.24e-01| 3.35e+00|Kkms |216|32| 1.01e+03| 1.57e+02| 5
IRASF17138-1017    |3| 2.62e+01| 1.32e+00| 3.94e+00|Kkms |185|22| 1.40e+03| 2.22e+02| 5
IRAS F17207-0014   |1| 7.00e+00| 0.00e+00| 1.40e+00|Kkms |   |44| 1.30e+02| 2.60e+01|12
IRAS F17207-0014   |1| 1.78e+02| 0.00e+00| 3.55e+01|Jykms|   |21| 1.99e+02| 3.99e+01| 7
IRAS F17207-0014   |1| 1.60e+02| 1.60e+01| 2.40e+01|Jykms|   |  |         |         |18
IRAS F17207-0014   |2| 3.27e+02| 3.70e+00| 6.54e+01|Jykms|   |13| 4.02e+02| 8.06e+01| 7
IRAS F17207-0014   |2| 6.88e+02| 1.09e+02| 1.03e+02|Jykms|   |  |         |         |18
IRAS F17207-0014   |3| 2.46e+01| 1.40e+00| 7.38e+00|Kkms |386|22| 1.14e+03| 3.49e+02|11
IRAS F17207-0014   |3| 1.20e+03| 1.90e+02| 1.80e+02|Jykms|   |  |         |         |18
IRAS F17207-0014   |4| 2.31e+03| 6.54e+02| 4.62e+02|Jykms|   |11| 2.93e+03| 1.02e+03|18
IRAS F17207-0014   |6| 3.40e+02| 1.40e+02| 8.50e+01|Jykms|   | 8| 4.56e+02| 2.20e+02|18
UGC11041           |1| 8.60e+00| 0.00e+00| 2.15e+00|Kkms |202|45| 1.79e+02| 4.47e+01| 1
UGC11041           |1| 4.21e+01| 0.00e+00| 1.05e+01|Kkms | 90|24| 3.12e+02| 7.81e+01| 1
UGC11041           |2| 1.04e+01| 0.00e+00| 2.60e+00|Kkms |159|24| 3.09e+02| 7.71e+01| 1
UGC11041           |2| 4.25e+01| 0.00e+00| 1.06e+01|Kkms |107|12| 4.54e+02| 1.13e+02| 1
IRAS17578-0400     |1| 6.71e+00| 6.55e-01| 1.01e+00|Kkms |237|55| 2.01e+02| 3.60e+01| 8
IRAS17578-0400     |2| 8.78e+00| 4.34e-01| 1.32e+00|Kkms |283|32| 3.99e+02| 6.31e+01| 5
IRAS17578-0400     |3| 1.57e+01| 6.98e-01| 2.36e+00|Kkms |194|22| 8.36e+02| 1.31e+02| 5
NGC6621            |1| 4.10e+00| 0.00e+00| 8.20e-01|Kkms |136|55| 1.16e+02| 2.32e+01| 2
IC4687             |1| 5.70e+00| 0.00e+00| 1.43e+00|Kkms | 68|45| 1.18e+02| 2.95e+01| 1
IC4687             |1| 6.00e+00| 0.00e+00| 1.20e+00|Kkms |   |44| 1.20e+02| 2.39e+01|12
IC4687             |1| 1.47e+02| 0.00e+00| 2.94e+01|Jykms|   |45| 1.45e+02| 2.91e+01| 7
IC4687             |1| 8.20e+00| 0.00e+00| 9.00e-01|Kkms |   |44| 1.63e+02| 1.79e+01| 3
IC4687             |2| 1.56e+01| 0.00e+00| 3.90e+00|Kkms |299|24| 4.62e+02| 1.15e+02| 1
IRAS F18293-3413   |1| 3.26e+01| 0.00e+00| 6.52e+00|Kkms |   |44| 6.49e+02| 1.30e+02|12
IRAS F18293-3413   |1| 3.63e+01| 4.00e-01| 3.63e+00|Kkms |261|45| 7.52e+02| 7.57e+01|13
IRAS F18293-3413   |1| 6.86e+02| 7.60e+00| 1.37e+02|Jykms|   |  |         |         | 7
IRAS F18293-3413   |2| 6.96e+01| 1.00e+00| 6.96e+00|Kkms |278|24| 1.91e+03| 1.93e+02|13
IRAS F18293-3413   |2| 1.43e+03| 2.05e+01| 2.85e+02|Jykms|   |  |         |         | 7
IC4734             |1| 1.16e+01| 0.00e+00| 2.32e+00|Kkms |   |44| 2.32e+02| 4.65e+01|12
IC4734             |1| 2.57e+02| 3.80e+00| 5.14e+01|Jykms|   |45| 2.55e+02| 5.11e+01| 7
IC4734             |1| 1.31e+01| 0.00e+00| 8.00e-01|Kkms |   |44| 2.62e+02| 1.60e+01| 3
IC4734             |1| 1.36e+01| 2.00e-01| 1.36e+00|Kkms |253|45| 2.83e+02| 2.86e+01|13
IC4734             |2| 1.50e+01| 6.00e-01| 1.50e+00|Kkms |217|24| 4.38e+02| 4.72e+01|13
IC4734             |2| 3.08e+02| 1.23e+01| 6.15e+01|Jykms|   |  |         |         | 7
NGC6701            |1| 6.70e+00| 0.00e+00| 1.34e+00|Kkms |100|55| 1.89e+02| 3.79e+01| 2
NGC6701            |1| 4.34e+01| 3.84e-01| 8.68e+00|Kkms |   |22| 3.31e+02| 6.63e+01| 4
NGC6701            |1| 3.81e+02| 0.00e+00| 7.62e+01|Jykms|   |22| 5.74e+02| 1.15e+02| 7
NGC6701            |1| 2.34e+02| 4.70e+01| 3.51e+01|Jykms|   |  |         |         |18
NGC6701            |2| 1.85e+01| 6.56e-01| 2.77e+00|Kkms |136|32| 9.35e+02| 1.44e+02| 5
NGC6701            |3| 2.26e+01| 1.60e+00| 3.39e+00|Kkms |122|22| 1.55e+03| 2.57e+02| 5
NGC6701            |3| 1.44e+03| 2.88e+02| 2.16e+02|Jykms|   |  |         |         |18
IRAS 19254-7245    |1| 2.40e+00| 0.00e+00| 4.80e-01|Kkms |   |44| 4.22e+01| 8.43e+00|12
IRAS 19254-7245    |1| 5.88e+01| 0.00e+00| 1.18e+01|Jykms|   |45| 5.84e+01| 1.17e+01| 7
IRAS 19297-0406    |3| 0.00e+00| 1.80e+00| 0.00e+00|Kkms |   |14| 0.00e+00| 4.86e+01|21
3C 405             |1| 0.00e+00| 1.90e+00| 0.00e+00|Jykms|   |55| 0.00e+00| 1.90e+00|19
MCG+04-48-002a     |1| 3.97e+00| 5.84e-01| 5.96e-01|Kkms |299|55| 1.17e+02| 2.46e+01| 8
MCG+04-48-002a     |2| 1.19e+01| 2.95e-01| 1.78e+00|Kkms |360|32| 5.51e+02| 8.38e+01| 5
MCG+04-48-002a     |3| 2.20e+01| 1.22e+00| 3.30e+00|Kkms |297|22| 1.23e+03| 1.97e+02| 5
NGC6946            |1| 1.43e+03| 0.00e+00| 2.86e+02|Jykms|   |22| 2.48e+03| 4.96e+02| 7
NGC6946            |2| 1.05e+02| 2.80e+00| 1.05e+01|Kkms |   |30| 5.63e+03| 5.83e+02|10
NGC6946            |3| 1.13e+02| 2.80e+00| 1.13e+01|Kkms |   |21| 9.25e+03| 9.53e+02|10
NGC6946            |3| 1.32e+02| 1.80e+00| 3.97e+01|Kkms |150|22| 1.09e+04| 3.26e+03|11
NGC6946            |4| 1.94e+02| 5.70e+00| 1.94e+01|Kkms |   |14| 1.74e+04| 1.82e+03|10
NGC6946            |6| 9.07e+01| 9.80e+00| 9.07e+00|Kkms |   |10| 1.27e+04| 1.87e+03|10
NGC6946_05         |2| 8.30e+00| 1.70e+00| 8.30e-01|Kkms |   |30| 5.08e+02| 1.16e+02|10
NGC6946_05         |3| 9.00e+00| 1.60e+00| 9.00e-01|Kkms |   |21| 9.60e+02| 1.96e+02|10
NGC6946_05         |4| 1.44e+01| 2.30e+00| 1.44e+00|Kkms |   |14| 2.16e+03| 4.07e+02|10
CGCG448-020        |1| 1.08e+01| 3.84e-01| 2.15e+00|Kkms |   |22| 6.60e+01| 1.34e+01| 4
CGCG448-020        |1| 8.03e+01| 0.00e+00| 1.61e+01|Jykms|   |21| 1.06e+02| 2.13e+01| 7
CGCG448-020        |1| 1.21e+02| 2.40e+01| 1.81e+01|Jykms|   |  |         |         |18
CGCG448-020        |2| 1.12e+02| 4.10e+00| 2.24e+01|Jykms|   |13| 1.91e+02| 3.88e+01| 7
CGCG448-020        |2| 7.25e+00| 4.88e-01| 1.09e+00|Kkms |190|32| 3.20e+02| 5.27e+01| 5
CGCG448-020        |3| 1.79e+01| 0.00e+00| 3.58e+00|Kkms |180|14| 5.06e+02| 1.01e+02|21
CGCG448-020        |3| 5.27e+02| 1.05e+02| 7.90e+01|Jykms|   |  |         |         |18
ESO286-IG019       |1| 3.10e+00| 0.00e+00| 6.20e-01|Kkms |   |44| 5.75e+01| 1.15e+01|12
3C 433             |1| 0.00e+00| 3.90e+00| 0.00e+00|Jykms|   |55| 0.00e+00| 3.90e+00|19
NGC7130            |1| 1.29e+01| 7.14e-01| 1.29e+00|Kkms |   |34| 1.67e+02| 1.90e+01|20
NGC7130            |1| 2.56e+02| 1.35e+01| 5.13e+01|Jykms|   |45| 2.54e+02| 5.25e+01| 7
NGC7130            |1| 9.35e+00| 5.20e-01| 9.35e-01|Kkms | 80|55| 2.73e+02| 3.12e+01| 6
NGC7130            |1| 1.43e+01| 0.00e+00| 5.00e-01|Kkms |   |44| 2.86e+02| 1.00e+01| 3
NGC7130            |1| 1.47e+01| 0.00e+00| 3.67e+00|Kkms | 85|45| 3.06e+02| 7.64e+01| 1
NGC7130            |2| 1.91e+01| 0.00e+00| 4.78e+00|Kkms | 96|24| 5.63e+02| 1.41e+02| 1
NGC7172            |1| 6.69e+00| 6.00e-01| 6.69e-01|Kkms |580|55| 1.94e+02| 2.60e+01| 6
NGC7172            |1| 1.58e+01| 0.00e+00| 3.95e+00|Kkms |216|45| 3.34e+02| 8.36e+01| 1
NGC7172            |2| 1.11e+01| 0.00e+00| 2.77e+00|Kkms |127|24| 3.52e+02| 8.80e+01| 1
ESO467-G027        |1| 7.10e+00| 0.00e+00| 1.77e+00|Kkms |132|45| 1.46e+02| 3.65e+01| 1
IC5179             |1| 2.87e+02| 5.70e+00| 5.75e+01|Jykms|   |45| 2.81e+02| 5.65e+01| 7
IC5179             |1| 1.40e+01| 0.00e+00| 2.80e+00|Kkms |   |44| 2.83e+02| 5.66e+01|12
IC5179             |1| 1.49e+01| 0.00e+00| 1.00e+00|Kkms |   |44| 3.01e+02| 2.02e+01| 3
IC5179             |1| 1.52e+01| 3.00e-01| 1.52e+00|Kkms |245|45| 3.17e+02| 3.23e+01|13
IC5179             |1| 2.02e+01| 0.00e+00| 5.05e+00|Kkms |166|45| 4.21e+02| 1.05e+02| 1
IC5179             |2| 4.02e+02| 1.23e+01| 8.04e+01|Jykms|   |24| 6.13e+02| 1.24e+02| 7
IC5179             |2| 1.96e+01| 6.00e-01| 1.96e+00|Kkms |209|24| 7.24e+02| 7.57e+01|13
IC5179             |2| 5.09e+01| 0.00e+00| 1.27e+01|Kkms |216|24| 1.88e+03| 4.70e+02| 1
NGC7331            |1| 2.69e+01| 0.00e+00| 3.70e+00|Kkms |   |33| 5.12e+02| 7.04e+01| 3
NGC7331            |1| 0.00e+00| 1.92e+02| 0.00e+00|Jykms|   |  |         |         | 7
NGC7331            |3| 7.20e+00| 6.00e-01| 2.16e+00|Kkms | 50|22| 1.24e+03| 3.85e+02|11
UGC12150           |1| 4.59e+00| 3.18e-01| 6.88e-01|Kkms |276|55| 1.34e+02| 2.22e+01| 8
UGC12150           |2| 1.23e+01| 5.92e-01| 1.85e+00|Kkms |309|32| 5.51e+02| 8.68e+01| 5
UGC12150           |3| 1.30e+01| 9.96e-01| 1.95e+00|Kkms |261|22| 6.83e+02| 1.15e+02| 5
IRAS 22491-1808    |1| 9.00e-01| 0.00e+00| 1.80e-01|Kkms |   |44| 1.52e+01| 3.03e+00|12
IRAS 22491-1808    |1| 2.20e+01| 0.00e+00| 4.40e+00|Jykms|   |45| 2.20e+01| 4.40e+00| 7
IRAS 22491-1808    |1| 9.00e-01| 0.00e+00| 1.80e-01|Kkms |135|55| 2.37e+01| 4.74e+00| 2
IRAS 22491-1808    |1| 3.30e+01| 6.00e+00| 4.95e+00|Jykms|   |  | 3.30e+01| 7.78e+00|18
IRAS 22491-1808    |2| 1.45e+02| 3.40e+01| 2.18e+01|Jykms|   |  | 1.45e+02| 4.04e+01|18
IRAS 22491-1808    |3| 5.58e+02| 1.90e+02| 8.37e+01|Jykms|   |  | 5.58e+02| 2.08e+02|18
NGC7465            |1| 1.19e+01| 4.46e-01| 2.38e+00|Kkms |   |21| 8.24e+01| 1.68e+01|24
NGC7465            |1| 5.30e+00| 2.90e-01| 5.30e-01|Kkms |110|55| 1.54e+02| 1.76e+01| 6
NGC7465            |2| 2.13e+01| 4.78e-01| 4.26e+00|Kkms |   |10| 2.11e+02| 4.25e+01|24
NGC7465            |3| 6.30e+00| 9.00e-01| 1.89e+00|Kkms |127|22| 4.04e+02| 1.34e+02|11
NGC7469            |1| 1.69e+01| 0.00e+00| 2.50e+00|Kkms |   |33| 2.06e+02| 3.05e+01| 3
NGC7469            |1| 9.60e+00| 0.00e+00| 1.92e+00|Kkms |200|55| 2.80e+02| 5.61e+01| 2
NGC7469            |1| 1.15e+01| 4.70e-01| 1.15e+00|Kkms |270|55| 3.36e+02| 3.63e+01| 6
NGC7469            |1| 2.98e+02| 2.70e+01| 4.47e+01|Jykms|   |  |         |         |18
NGC7469            |1| 4.81e+01| 0.00e+00| 9.62e+00|Jykms|   |  |         |         | 7
NGC7469            |2| 5.92e+01| 2.03e+00| 8.89e+00|Kkms |257|32| 2.75e+03| 4.23e+02| 5
NGC7469            |2| 8.90e+02| 1.03e+02| 1.34e+02|Jykms|   |  |         |         |18
NGC7469            |3| 3.52e+01| 1.30e+00| 1.06e+01|Kkms |249|22| 1.98e+03| 5.99e+02|11
NGC7469            |3| 1.60e+03| 2.40e+02| 2.40e+02|Jykms|   |  |         |         |18
NGC7469            |4| 3.97e+03| 8.20e+02| 7.94e+02|Jykms|   |11| 6.55e+03| 1.88e+03|18
NGC7469            |6| 2.36e+03| 5.90e+02| 5.89e+02|Jykms|   | 8| 4.40e+03| 1.56e+03|18
ESO148-IG002       |1| 1.90e+00| 0.00e+00| 3.80e-01|Kkms |   |44| 3.50e+01| 7.01e+00|12
ESO148-IG002       |1| 4.65e+01| 0.00e+00| 9.30e+00|Jykms|   |45| 4.62e+01| 9.24e+00| 7
IC5298             |1| 2.40e+00| 0.00e+00| 4.80e-01|Kkms |214|55| 6.95e+01| 1.39e+01| 2
IC5298             |2| 3.97e+00| 1.74e-01| 5.95e-01|Kkms |261|32| 1.72e+02| 2.68e+01| 5
IC5298             |3| 4.86e+00| 5.26e-01| 7.30e-01|Kkms |179|22| 2.40e+02| 4.44e+01| 5
NGC7552            |1| 4.00e+01| 7.14e-01| 4.00e+00|Kkms |   |34| 5.43e+02| 5.51e+01|20
NGC7552            |1| 6.52e+02| 8.81e+01| 1.30e+02|Jykms|   |45| 6.44e+02| 1.55e+02| 7
NGC7552            |1| 4.19e+01| 8.00e-01| 4.19e+00|Kkms |305|45| 8.97e+02| 9.13e+01|40
NGC7552            |2| 1.23e+02| 1.60e+00| 1.23e+01|Kkms |   |24| 3.75e+03| 3.78e+02|20
NGC7591            |1| 2.96e+01| 3.72e-01| 5.92e+00|Kkms |   |22| 2.06e+02| 4.12e+01| 4
NGC7591            |2| 1.18e+01| 5.60e-01| 1.78e+00|Kkms |354|32| 5.78e+02| 9.08e+01| 5
NGC7591            |3| 3.93e+01| 7.24e-01| 5.90e+00|Kkms |309|22| 2.46e+03| 3.72e+02| 5
NGC7592            |1| 1.73e+01| 0.00e+00| 4.33e+00|Kkms |258|24| 1.30e+02| 3.24e+01| 1
NGC7592            |1| 5.90e+00| 0.00e+00| 1.18e+00|Kkms |259|55| 1.67e+02| 3.34e+01| 2
NGC7592            |2| 3.82e+01| 0.00e+00| 9.55e+00|Kkms |266|12| 4.66e+02| 1.17e+02| 1
NGC7592            |3| 0.00e+00| 6.20e+00| 0.00e+00|Kkms |   |14| 0.00e+00| 2.05e+02|21
NGC7582            |1| 3.00e+01| 1.43e+00| 3.00e+00|Kkms |   |34| 4.16e+02| 4.61e+01|20
NGC7582            |1| 6.96e+02| 6.90e+01| 1.39e+02|Jykms|   |45| 6.85e+02| 1.53e+02| 7
NGC7582            |1| 3.97e+01| 7.00e-01| 3.97e+00|Kkms |420|45| 8.47e+02| 8.60e+01|40
NGC7582            |2| 1.16e+02| 4.00e+00| 1.16e+01|Kkms |   |24| 3.81e+03| 4.04e+02|20
NGC7674            |1| 3.85e+00| 2.10e-01| 3.85e-01|Kkms |195|55| 1.03e+02| 1.18e+01| 6
NGC7674            |1| 4.00e+00| 0.00e+00| 8.00e-01|Kkms |145|55| 1.07e+02| 2.15e+01| 2
NGC7679a           |1| 3.36e+00| 2.66e-01| 5.03e-01|Kkms |184|55| 9.70e+01| 1.64e+01| 8
NGC7679a           |3| 1.72e+01| 1.40e+00| 5.16e+00|Kkms |285|22| 1.01e+03| 3.15e+02|11
IRAS 23365+3604    |1| 4.21e+01| 0.00e+00| 8.42e+00|Jykms|   |21| 4.62e+01| 9.23e+00| 7
IRAS 23365+3604    |1| 1.07e+01| 0.00e+00| 2.14e+00|Kkms |310|22| 5.09e+01| 1.02e+01|17
IRAS 23365+3604    |1| 3.90e+01| 6.00e+00| 5.85e+00|Jykms|   |  |         |         |18
IRAS 23365+3604    |2| 1.17e+02| 2.00e+01| 1.76e+01|Jykms|   |  |         |         |18
IRAS 23365+3604    |3| 2.88e+02| 7.10e+01| 4.32e+01|Jykms|   |  |         |         |18
IRAS 23365+3604    |4| 0.00e+00| 4.89e+02| 0.00e+00|Jykms|   |11| 0.00e+00| 5.77e+02|18
IRAS 23365+3604    |6| 2.95e+02| 1.10e+02| 7.38e+01|Jykms|   | 8| 3.59e+02| 1.61e+02|18
NGC7771            |1| 1.20e+01| 0.00e+00| 2.40e+00|Kkms |300|55| 3.42e+02| 6.84e+01| 2
NGC7771            |1| 3.12e+01| 0.00e+00| 2.10e+00|Kkms |   |33| 3.96e+02| 2.67e+01| 3
NGC7771            |1| 4.96e+02| 0.00e+00| 9.92e+01|Jykms|   |21| 6.58e+02| 1.32e+02| 7
NGC7771            |2| 4.16e+01| 4.34e-01| 6.24e+00|Kkms |343|32| 2.01e+03| 3.02e+02| 5
NGC7771            |3| 3.84e+01| 5.14e-01| 5.76e+00|Kkms |330|22| 2.27e+03| 3.43e+02| 5
Mrk331             |1| 4.95e+01| 0.00e+00| 9.90e+00|Jykms|   |21| 5.94e+01| 1.19e+01| 7
Mrk331             |1| 1.16e+01| 0.00e+00| 2.32e+00|Kkms |245|55| 3.42e+02| 6.84e+01| 2
Mrk331             |2| 1.28e+01| 4.52e-01| 1.92e+00|Kkms |290|32| 5.77e+02| 8.89e+01| 5
Mrk331             |3| 2.80e+01| 9.97e-01| 4.20e+00|Kkms |291|22| 1.49e+03| 2.29e+02| 5

